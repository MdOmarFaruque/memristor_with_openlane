VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO core_flat_v4
  CLASS BLOCK ;
  FOREIGN core_flat_v4 ;
  ORIGIN 400.150 350.900 ;
  SIZE 650.000 BY 679.000 ;
  PIN SEL1
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT -287.380 -15.150 -287.050 -14.980 ;
        RECT -255.700 -16.340 -255.370 -16.170 ;
        RECT -287.380 -16.700 -287.050 -16.530 ;
        RECT -255.700 -17.890 -255.370 -17.720 ;
        RECT -287.330 -18.470 -287.000 -18.300 ;
        RECT -287.330 -20.110 -287.000 -19.940 ;
        RECT -255.680 -19.980 -255.350 -19.810 ;
        RECT -255.680 -21.620 -255.350 -21.450 ;
      LAYER mcon ;
        RECT -287.300 -15.150 -287.130 -14.980 ;
        RECT -255.620 -16.340 -255.450 -16.170 ;
        RECT -287.300 -16.700 -287.130 -16.530 ;
        RECT -255.620 -17.890 -255.450 -17.720 ;
        RECT -287.250 -18.470 -287.080 -18.300 ;
        RECT -287.250 -20.110 -287.080 -19.940 ;
        RECT -255.600 -19.980 -255.430 -19.810 ;
        RECT -255.600 -21.620 -255.430 -21.450 ;
      LAYER met1 ;
        RECT -289.540 -8.750 -289.020 -8.660 ;
        RECT -276.860 -8.750 -273.060 -8.720 ;
        RECT -262.050 -8.750 -258.230 -7.530 ;
        RECT -289.650 -9.170 -258.230 -8.750 ;
        RECT -289.540 -13.020 -289.020 -9.170 ;
        RECT -262.050 -9.880 -258.230 -9.170 ;
        RECT -289.550 -13.220 -289.020 -13.020 ;
        RECT -298.220 -17.350 -296.360 -16.750 ;
        RECT -299.830 -17.460 -289.780 -17.350 ;
        RECT -289.550 -17.460 -289.030 -13.220 ;
        RECT -287.420 -15.190 -287.030 -14.890 ;
        RECT -262.120 -15.650 -258.700 -14.060 ;
        RECT -287.430 -17.430 -286.980 -16.500 ;
        RECT -288.580 -17.460 -286.980 -17.430 ;
        RECT -299.830 -17.680 -286.980 -17.460 ;
        RECT -299.830 -17.770 -289.780 -17.680 ;
        RECT -288.580 -17.690 -286.980 -17.680 ;
        RECT -298.220 -18.280 -296.360 -17.770 ;
        RECT -287.430 -18.510 -286.980 -17.690 ;
        RECT -287.370 -18.520 -286.980 -18.510 ;
        RECT -261.370 -18.490 -260.160 -15.650 ;
        RECT -259.620 -16.110 -257.910 -16.100 ;
        RECT -255.700 -16.110 -255.370 -16.070 ;
        RECT -259.620 -16.350 -255.370 -16.110 ;
        RECT -259.620 -18.490 -259.070 -16.350 ;
        RECT -258.410 -16.360 -255.370 -16.350 ;
        RECT -255.680 -16.370 -255.390 -16.360 ;
        RECT -255.700 -17.960 -255.370 -17.680 ;
        RECT -261.370 -19.030 -259.070 -18.490 ;
        RECT -260.850 -19.040 -259.070 -19.030 ;
        RECT -287.370 -20.150 -286.980 -19.880 ;
        RECT -259.620 -21.430 -259.070 -19.040 ;
        RECT -255.670 -20.000 -255.340 -19.720 ;
        RECT -255.660 -20.010 -255.370 -20.000 ;
        RECT -255.670 -21.430 -255.340 -21.400 ;
        RECT -259.620 -21.740 -255.330 -21.430 ;
        RECT -259.620 -21.750 -259.070 -21.740 ;
      LAYER via ;
        RECT -261.010 -8.860 -259.710 -8.190 ;
        RECT -297.690 -17.810 -297.140 -17.300 ;
        RECT -261.200 -14.990 -260.240 -14.600 ;
      LAYER met2 ;
        RECT -261.380 -9.640 -259.470 -7.710 ;
        RECT -261.380 -9.660 -260.160 -9.640 ;
        RECT -261.260 -14.200 -260.160 -9.660 ;
        RECT -259.950 -9.660 -259.470 -9.640 ;
        RECT -259.950 -9.680 -259.660 -9.660 ;
        RECT -261.280 -14.290 -260.160 -14.200 ;
        RECT -261.280 -15.540 -260.090 -14.290 ;
        RECT -300.590 -17.180 -299.350 -17.020 ;
        RECT -298.160 -17.180 -296.450 -16.920 ;
        RECT -300.590 -17.880 -296.450 -17.180 ;
        RECT -300.590 -18.220 -299.350 -17.880 ;
        RECT -298.160 -18.110 -296.450 -17.880 ;
      LAYER via2 ;
        RECT -300.260 -17.880 -299.770 -17.450 ;
      LAYER met3 ;
        RECT -392.160 -17.190 -390.160 -17.180 ;
        RECT -300.430 -17.190 -299.540 -17.180 ;
        RECT -392.160 -17.780 -299.540 -17.190 ;
        RECT -300.430 -18.070 -299.540 -17.780 ;
    END
  END SEL1
  PIN DIGITALIN1
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT -272.530 -16.070 -272.200 -15.900 ;
        RECT -252.240 -16.230 -251.910 -16.060 ;
        RECT -272.530 -17.620 -272.200 -17.450 ;
        RECT -252.240 -17.780 -251.910 -17.610 ;
        RECT -272.550 -19.840 -272.220 -19.670 ;
        RECT -252.260 -20.000 -251.930 -19.830 ;
        RECT -272.550 -21.480 -272.220 -21.310 ;
        RECT -252.260 -21.640 -251.930 -21.470 ;
      LAYER mcon ;
        RECT -272.450 -16.070 -272.280 -15.900 ;
        RECT -252.160 -16.230 -251.990 -16.060 ;
        RECT -272.450 -17.620 -272.280 -17.450 ;
        RECT -252.160 -17.780 -251.990 -17.610 ;
        RECT -272.470 -19.840 -272.300 -19.670 ;
        RECT -252.180 -20.000 -252.010 -19.830 ;
        RECT -272.470 -21.480 -272.300 -21.310 ;
        RECT -252.180 -21.640 -252.010 -21.470 ;
      LAYER met1 ;
        RECT -272.530 -16.110 -272.200 -15.830 ;
        RECT -252.240 -16.270 -251.910 -15.990 ;
        RECT -270.300 -17.410 -269.700 -17.390 ;
        RECT -272.540 -17.680 -269.700 -17.410 ;
        RECT -250.010 -17.570 -249.410 -17.550 ;
        RECT -272.540 -17.690 -269.740 -17.680 ;
        RECT -272.550 -19.870 -272.220 -19.590 ;
        RECT -270.240 -21.280 -269.740 -17.690 ;
        RECT -252.250 -17.840 -249.410 -17.570 ;
        RECT -252.250 -17.850 -249.450 -17.840 ;
        RECT -252.260 -20.030 -251.930 -19.750 ;
        RECT -272.580 -21.630 -269.740 -21.280 ;
        RECT -249.950 -21.440 -249.450 -17.850 ;
        RECT -270.240 -22.080 -269.740 -21.630 ;
        RECT -252.290 -21.790 -249.450 -21.440 ;
        RECT -270.210 -22.450 -269.760 -22.080 ;
        RECT -249.950 -22.240 -249.450 -21.790 ;
        RECT -270.520 -23.030 -269.560 -22.450 ;
        RECT -249.920 -22.610 -249.470 -22.240 ;
        RECT -250.230 -23.190 -249.270 -22.610 ;
        RECT -270.790 -24.320 -269.550 -24.120 ;
        RECT -270.830 -25.540 -267.840 -24.320 ;
        RECT -250.500 -24.410 -249.260 -24.280 ;
        RECT -250.790 -25.750 -248.300 -24.410 ;
        RECT -260.850 -34.320 -258.060 -32.950 ;
        RECT -261.140 -37.020 -257.780 -34.320 ;
      LAYER via ;
        RECT -270.300 -22.880 -269.870 -22.620 ;
        RECT -250.010 -23.040 -249.580 -22.780 ;
        RECT -270.460 -24.650 -270.020 -24.390 ;
        RECT -270.360 -25.110 -268.760 -24.720 ;
        RECT -250.170 -24.810 -249.730 -24.550 ;
        RECT -250.270 -25.180 -249.230 -24.920 ;
        RECT -260.450 -33.990 -258.740 -33.430 ;
        RECT -259.930 -36.100 -258.910 -35.440 ;
      LAYER met2 ;
        RECT -299.490 -19.060 -298.460 -18.990 ;
        RECT -299.490 -19.680 -294.420 -19.060 ;
        RECT -299.490 -19.940 -298.460 -19.680 ;
        RECT -295.270 -35.320 -294.420 -19.680 ;
        RECT -270.430 -22.950 -269.660 -22.530 ;
        RECT -270.370 -24.210 -269.800 -22.950 ;
        RECT -250.140 -23.110 -249.370 -22.690 ;
        RECT -270.700 -24.520 -269.630 -24.210 ;
        RECT -250.080 -24.370 -249.510 -23.110 ;
        RECT -270.700 -24.840 -268.020 -24.520 ;
        RECT -250.410 -24.580 -249.340 -24.370 ;
        RECT -270.680 -25.430 -268.020 -24.840 ;
        RECT -270.420 -27.040 -268.630 -25.430 ;
        RECT -250.630 -25.520 -248.610 -24.580 ;
        RECT -250.230 -27.040 -248.960 -25.520 ;
        RECT -270.540 -27.280 -248.960 -27.040 ;
        RECT -270.540 -27.300 -249.540 -27.280 ;
        RECT -260.190 -27.320 -258.480 -27.300 ;
        RECT -260.190 -33.130 -259.380 -27.320 ;
        RECT -260.680 -33.140 -259.380 -33.130 ;
        RECT -260.680 -33.170 -258.700 -33.140 ;
        RECT -260.680 -34.370 -258.220 -33.170 ;
        RECT -260.880 -35.270 -257.940 -34.780 ;
        RECT -272.670 -35.320 -257.940 -35.270 ;
        RECT -295.270 -36.160 -257.940 -35.320 ;
        RECT -295.270 -36.210 -272.550 -36.160 ;
        RECT -295.270 -36.330 -294.420 -36.210 ;
        RECT -260.880 -36.860 -257.940 -36.160 ;
      LAYER via2 ;
        RECT -299.300 -19.730 -298.720 -19.200 ;
      LAYER met3 ;
        RECT -299.390 -19.250 -298.580 -19.080 ;
        RECT -392.130 -19.840 -298.580 -19.250 ;
        RECT -392.130 -19.850 -390.130 -19.840 ;
        RECT -299.390 -19.870 -298.580 -19.840 ;
    END
  END DIGITALIN1
  PIN AIN1
    ANTENNADIFFAREA 23.199999 ;
    PORT
      LAYER li1 ;
        RECT -162.830 7.935 -162.660 27.975 ;
        RECT -158.390 8.130 -158.220 28.170 ;
        RECT -164.120 -58.625 -163.950 -38.585 ;
        RECT -159.680 -58.430 -159.510 -38.390 ;
      LAYER mcon ;
        RECT -162.830 8.015 -162.660 27.895 ;
        RECT -158.390 8.210 -158.220 28.090 ;
        RECT -164.120 -58.545 -163.950 -38.665 ;
        RECT -159.680 -58.350 -159.510 -38.470 ;
      LAYER met1 ;
        RECT -162.860 8.910 -162.630 27.955 ;
        RECT -164.740 8.900 -162.630 8.910 ;
        RECT -165.510 8.750 -162.630 8.900 ;
        RECT -168.020 8.700 -162.630 8.750 ;
        RECT -168.090 8.350 -162.630 8.700 ;
        RECT -168.090 -8.270 -167.740 8.350 ;
        RECT -165.510 8.000 -162.630 8.350 ;
        RECT -158.420 8.590 -158.190 28.150 ;
        RECT -157.130 8.590 -156.270 8.700 ;
        RECT -158.420 8.240 -156.270 8.590 ;
        RECT -158.420 8.150 -158.190 8.240 ;
        RECT -165.510 7.990 -163.400 8.000 ;
        RECT -165.130 5.640 -164.420 7.990 ;
        RECT -162.860 7.955 -162.630 8.000 ;
        RECT -157.130 5.640 -156.270 8.240 ;
        RECT -165.130 5.070 -156.270 5.640 ;
        RECT -165.130 4.960 -156.280 5.070 ;
        RECT -165.110 4.950 -156.280 4.960 ;
        RECT -150.340 -8.270 -144.570 -5.490 ;
        RECT -168.090 -9.660 -144.570 -8.270 ;
        RECT -168.090 -35.710 -167.740 -9.660 ;
        RECT -150.340 -12.670 -144.570 -9.660 ;
        RECT -168.840 -36.900 -166.930 -35.710 ;
        RECT -169.060 -48.290 -167.260 -46.930 ;
        RECT -168.790 -58.220 -167.910 -48.290 ;
        RECT -164.150 -57.650 -163.920 -38.605 ;
        RECT -166.030 -57.660 -163.920 -57.650 ;
        RECT -166.800 -58.220 -163.920 -57.660 ;
        RECT -168.860 -58.560 -163.920 -58.220 ;
        RECT -159.710 -57.970 -159.480 -38.410 ;
        RECT -158.420 -57.970 -157.560 -57.860 ;
        RECT -159.710 -58.320 -157.560 -57.970 ;
        RECT -159.710 -58.410 -159.480 -58.320 ;
        RECT -168.860 -58.570 -164.690 -58.560 ;
        RECT -166.420 -60.920 -165.710 -58.570 ;
        RECT -164.150 -58.605 -163.920 -58.560 ;
        RECT -158.420 -60.920 -157.560 -58.320 ;
        RECT -166.420 -61.490 -157.560 -60.920 ;
        RECT -166.420 -61.600 -157.570 -61.490 ;
        RECT -166.400 -61.610 -157.570 -61.600 ;
      LAYER via ;
        RECT -148.560 -9.740 -146.640 -8.420 ;
        RECT -168.400 -36.460 -167.880 -36.120 ;
        RECT -168.580 -47.730 -168.010 -47.430 ;
      LAYER met2 ;
        RECT -284.210 92.620 -132.160 92.970 ;
        RECT -284.390 91.380 -132.160 92.620 ;
        RECT -284.390 0.780 -282.980 91.380 ;
        RECT -299.480 -0.020 -282.830 0.780 ;
        RECT -301.360 -12.320 -299.820 -12.180 ;
        RECT -299.480 -12.320 -298.730 -0.020 ;
        RECT -149.730 -7.990 -145.180 -6.190 ;
        RECT -134.620 -7.990 -132.660 91.380 ;
        RECT -149.730 -9.950 -132.660 -7.990 ;
        RECT -149.730 -11.880 -145.180 -9.950 ;
        RECT -134.620 -10.740 -132.660 -9.950 ;
        RECT -301.360 -13.390 -298.640 -12.320 ;
        RECT -301.360 -13.590 -299.820 -13.390 ;
        RECT -299.480 -13.430 -298.730 -13.390 ;
        RECT -168.760 -36.770 -167.120 -35.820 ;
        RECT -168.520 -47.000 -167.690 -36.770 ;
        RECT -168.990 -48.230 -167.400 -47.000 ;
      LAYER via2 ;
        RECT -301.070 -13.280 -300.310 -12.550 ;
      LAYER met3 ;
        RECT -392.160 -12.480 -390.140 -12.470 ;
        RECT -301.200 -12.480 -299.960 -12.340 ;
        RECT -392.160 -13.070 -299.770 -12.480 ;
        RECT -301.200 -13.470 -299.960 -13.070 ;
    END
  END AIN1
  PIN SEL3
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT 45.430 -205.420 45.600 -205.090 ;
        RECT 46.980 -205.420 47.150 -205.090 ;
        RECT 49.070 -205.400 49.240 -205.070 ;
        RECT 50.710 -205.400 50.880 -205.070 ;
        RECT 44.240 -237.100 44.410 -236.770 ;
        RECT 45.790 -237.100 45.960 -236.770 ;
        RECT 47.560 -237.050 47.730 -236.720 ;
        RECT 49.200 -237.050 49.370 -236.720 ;
      LAYER mcon ;
        RECT 45.430 -205.340 45.600 -205.170 ;
        RECT 46.980 -205.340 47.150 -205.170 ;
        RECT 49.070 -205.320 49.240 -205.150 ;
        RECT 50.710 -205.320 50.880 -205.150 ;
        RECT 44.240 -237.020 44.410 -236.850 ;
        RECT 45.790 -237.020 45.960 -236.850 ;
        RECT 47.560 -236.970 47.730 -236.800 ;
        RECT 49.200 -236.970 49.370 -236.800 ;
      LAYER met1 ;
        RECT 50.690 -205.060 51.000 -205.050 ;
        RECT 48.980 -205.090 49.260 -205.060 ;
        RECT 45.330 -205.110 45.620 -205.090 ;
        RECT 45.330 -205.400 45.630 -205.110 ;
        RECT 45.330 -205.420 45.620 -205.400 ;
        RECT 46.940 -205.420 47.220 -205.090 ;
        RECT 48.980 -205.380 49.270 -205.090 ;
        RECT 48.980 -205.390 49.260 -205.380 ;
        RECT 50.660 -205.390 51.000 -205.060 ;
        RECT 45.370 -207.630 45.620 -205.420 ;
        RECT 36.790 -211.770 39.140 -207.950 ;
        RECT 45.360 -208.130 45.620 -207.630 ;
        RECT 43.320 -209.880 44.910 -208.420 ;
        RECT 45.360 -208.790 45.610 -208.130 ;
        RECT 50.690 -208.790 51.000 -205.390 ;
        RECT 45.360 -209.340 51.010 -208.790 ;
        RECT 47.750 -209.880 48.300 -209.340 ;
        RECT 43.320 -210.570 48.300 -209.880 ;
        RECT 43.320 -211.090 48.290 -210.570 ;
        RECT 38.010 -222.780 38.430 -211.770 ;
        RECT 43.320 -211.840 44.910 -211.090 ;
        RECT 37.980 -226.580 38.430 -222.780 ;
        RECT 38.010 -238.740 38.430 -226.580 ;
        RECT 44.150 -237.140 44.450 -236.750 ;
        RECT 45.760 -237.090 47.780 -236.700 ;
        RECT 49.140 -237.090 49.410 -236.700 ;
        RECT 45.760 -237.150 47.770 -237.090 ;
        RECT 46.690 -238.300 46.950 -237.150 ;
        RECT 37.920 -238.750 42.480 -238.740 ;
        RECT 46.720 -238.750 46.940 -238.300 ;
        RECT 37.920 -239.260 46.940 -238.750 ;
        RECT 38.010 -239.370 38.430 -239.260 ;
        RECT 42.280 -239.270 46.940 -239.260 ;
        RECT 46.720 -239.500 46.940 -239.270 ;
        RECT 46.610 -248.990 47.030 -239.500 ;
        RECT 46.370 -249.950 47.310 -248.990 ;
      LAYER via ;
        RECT 37.450 -210.730 38.120 -209.430 ;
        RECT 43.860 -210.920 44.250 -209.960 ;
        RECT 46.720 -249.620 46.980 -249.360 ;
      LAYER met2 ;
        RECT 36.970 -209.380 38.920 -209.190 ;
        RECT 36.970 -209.670 38.940 -209.380 ;
        RECT 36.970 -209.880 38.900 -209.670 ;
        RECT 43.550 -209.880 44.800 -209.810 ;
        RECT 36.970 -210.980 44.800 -209.880 ;
        RECT 36.970 -211.100 38.920 -210.980 ;
        RECT 43.460 -211.000 44.800 -210.980 ;
        RECT 46.240 -348.890 47.590 -248.940 ;
        RECT 46.690 -350.900 46.990 -348.890 ;
    END
  END SEL3
  PIN DIGITALIN3
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT 45.320 -201.960 45.490 -201.630 ;
        RECT 46.870 -201.960 47.040 -201.630 ;
        RECT 49.090 -201.980 49.260 -201.650 ;
        RECT 50.730 -201.980 50.900 -201.650 ;
        RECT 45.160 -222.250 45.330 -221.920 ;
        RECT 46.710 -222.250 46.880 -221.920 ;
        RECT 48.930 -222.270 49.100 -221.940 ;
        RECT 50.570 -222.270 50.740 -221.940 ;
      LAYER mcon ;
        RECT 45.320 -201.880 45.490 -201.710 ;
        RECT 46.870 -201.880 47.040 -201.710 ;
        RECT 49.090 -201.900 49.260 -201.730 ;
        RECT 50.730 -201.900 50.900 -201.730 ;
        RECT 45.160 -222.170 45.330 -222.000 ;
        RECT 46.710 -222.170 46.880 -222.000 ;
        RECT 48.930 -222.190 49.100 -222.020 ;
        RECT 50.570 -222.190 50.740 -222.020 ;
      LAYER met1 ;
        RECT 53.670 -198.980 55.010 -198.020 ;
        RECT 46.810 -199.170 47.100 -199.130 ;
        RECT 46.810 -199.190 51.500 -199.170 ;
        RECT 51.870 -199.190 52.450 -198.990 ;
        RECT 46.810 -199.640 52.450 -199.190 ;
        RECT 46.810 -199.670 51.500 -199.640 ;
        RECT 46.810 -199.730 47.110 -199.670 ;
        RECT 45.250 -201.960 45.530 -201.630 ;
        RECT 46.830 -201.970 47.110 -199.730 ;
        RECT 49.010 -201.980 49.290 -201.650 ;
        RECT 50.700 -202.010 51.050 -199.670 ;
        RECT 51.870 -199.950 52.450 -199.640 ;
        RECT 53.540 -200.220 55.010 -198.980 ;
        RECT 53.670 -200.510 55.010 -200.220 ;
        RECT 63.580 -207.780 66.280 -207.500 ;
        RECT 62.210 -210.570 66.280 -207.780 ;
        RECT 63.580 -210.860 66.280 -210.570 ;
        RECT 53.580 -219.270 54.800 -217.560 ;
        RECT 46.650 -219.460 46.940 -219.420 ;
        RECT 46.650 -219.480 51.340 -219.460 ;
        RECT 51.710 -219.480 52.290 -219.280 ;
        RECT 46.650 -219.930 52.290 -219.480 ;
        RECT 46.650 -219.960 51.340 -219.930 ;
        RECT 46.650 -220.020 46.950 -219.960 ;
        RECT 45.090 -222.250 45.370 -221.920 ;
        RECT 46.670 -222.260 46.950 -220.020 ;
        RECT 48.850 -222.270 49.130 -221.940 ;
        RECT 50.540 -222.300 50.890 -219.960 ;
        RECT 51.710 -220.240 52.290 -219.930 ;
        RECT 53.380 -220.510 54.800 -219.270 ;
        RECT 53.580 -220.550 54.800 -220.510 ;
      LAYER via ;
        RECT 52.040 -199.730 52.300 -199.300 ;
        RECT 53.810 -199.890 54.070 -199.450 ;
        RECT 54.180 -199.990 54.440 -198.950 ;
        RECT 62.690 -210.170 63.250 -208.460 ;
        RECT 64.700 -209.650 65.360 -208.630 ;
        RECT 51.880 -220.020 52.140 -219.590 ;
        RECT 53.650 -220.180 53.910 -219.740 ;
        RECT 53.980 -220.080 54.370 -218.480 ;
      LAYER met2 ;
        RECT 53.840 -198.680 54.780 -198.330 ;
        RECT 53.840 -199.060 56.540 -198.680 ;
        RECT 51.950 -199.230 52.370 -199.090 ;
        RECT 53.630 -199.230 56.540 -199.060 ;
        RECT 51.950 -199.260 56.540 -199.230 ;
        RECT 51.950 -199.800 56.560 -199.260 ;
        RECT 51.950 -199.860 52.370 -199.800 ;
        RECT 53.630 -199.950 56.560 -199.800 ;
        RECT 53.630 -200.130 54.780 -199.950 ;
        RECT 53.840 -200.350 54.780 -200.130 ;
        RECT 56.300 -208.200 56.560 -199.950 ;
        RECT 56.300 -209.100 56.580 -208.200 ;
        RECT 62.430 -208.420 63.630 -207.940 ;
        RECT 62.400 -209.100 63.630 -208.420 ;
        RECT 56.300 -209.910 63.630 -209.100 ;
        RECT 53.780 -218.350 54.690 -217.740 ;
        RECT 56.300 -218.350 56.560 -209.910 ;
        RECT 62.390 -210.400 63.630 -209.910 ;
        RECT 64.040 -210.600 66.120 -207.660 ;
        RECT 53.780 -219.350 56.560 -218.350 ;
        RECT 51.790 -219.520 52.210 -219.380 ;
        RECT 53.470 -219.520 56.560 -219.350 ;
        RECT 51.790 -220.090 56.560 -219.520 ;
        RECT 51.790 -220.150 52.210 -220.090 ;
        RECT 53.470 -220.140 56.560 -220.090 ;
        RECT 53.470 -220.400 54.690 -220.140 ;
        RECT 56.300 -220.260 56.560 -220.140 ;
        RECT 53.470 -220.420 54.100 -220.400 ;
        RECT 64.530 -222.270 65.420 -210.600 ;
        RECT 64.530 -222.390 65.470 -222.270 ;
        RECT 64.580 -244.140 65.470 -222.390 ;
        RECT 48.320 -244.990 65.590 -244.140 ;
        RECT 48.320 -248.090 48.940 -244.990 ;
        RECT 49.650 -248.090 51.100 -248.050 ;
        RECT 48.310 -248.660 51.100 -248.090 ;
        RECT 49.650 -249.070 51.100 -248.660 ;
        RECT 49.690 -348.890 51.040 -249.070 ;
        RECT 50.250 -350.890 50.550 -348.890 ;
    END
  END DIGITALIN3
  PIN AIN3
    ANTENNADIFFAREA 23.199999 ;
    PORT
      LAYER li1 ;
        RECT 1.090 -108.110 21.130 -107.940 ;
        RECT 67.650 -109.400 87.690 -109.230 ;
        RECT 1.285 -112.550 21.325 -112.380 ;
        RECT 67.845 -113.840 87.885 -113.670 ;
      LAYER mcon ;
        RECT 1.170 -108.110 21.050 -107.940 ;
        RECT 67.730 -109.400 87.610 -109.230 ;
        RECT 1.365 -112.550 21.245 -112.380 ;
        RECT 67.925 -113.840 87.805 -113.670 ;
      LAYER met1 ;
        RECT 34.750 -100.060 41.930 -94.290 ;
        RECT 20.560 -106.000 24.190 -105.990 ;
        RECT 20.560 -106.850 24.310 -106.000 ;
        RECT 20.670 -107.910 21.020 -106.850 ;
        RECT 1.110 -108.140 21.110 -107.910 ;
        RECT 1.305 -112.580 21.305 -112.350 ;
        RECT 20.350 -113.120 21.260 -112.580 ;
        RECT 20.350 -114.140 21.270 -113.120 ;
        RECT 23.620 -114.140 24.310 -106.850 ;
        RECT 20.350 -114.460 24.310 -114.140 ;
        RECT 20.360 -114.830 24.310 -114.460 ;
        RECT 20.360 -114.850 24.300 -114.830 ;
        RECT 20.360 -115.230 21.270 -114.850 ;
        RECT 20.510 -117.460 20.910 -115.230 ;
        RECT 37.530 -117.460 38.920 -100.060 ;
        RECT 87.120 -107.290 90.750 -107.280 ;
        RECT 87.120 -108.140 90.870 -107.290 ;
        RECT 87.230 -109.200 87.580 -108.140 ;
        RECT 67.670 -109.430 87.670 -109.200 ;
        RECT 67.865 -113.870 87.865 -113.640 ;
        RECT 86.910 -114.410 87.820 -113.870 ;
        RECT 86.910 -115.430 87.830 -114.410 ;
        RECT 90.180 -115.430 90.870 -108.140 ;
        RECT 86.910 -115.750 90.870 -115.430 ;
        RECT 86.920 -116.120 90.870 -115.750 ;
        RECT 86.920 -116.140 90.860 -116.120 ;
        RECT 86.920 -116.520 87.830 -116.140 ;
        RECT 64.970 -117.460 66.160 -116.650 ;
        RECT 20.510 -117.740 66.160 -117.460 ;
        RECT 20.560 -117.810 66.160 -117.740 ;
        RECT 64.970 -118.560 66.160 -117.810 ;
        RECT 76.190 -117.630 77.550 -116.980 ;
        RECT 87.480 -117.630 87.830 -116.520 ;
        RECT 76.190 -118.510 87.830 -117.630 ;
        RECT 76.190 -118.780 77.550 -118.510 ;
        RECT 87.480 -118.580 87.830 -118.510 ;
      LAYER via ;
        RECT 37.680 -98.280 39.000 -96.360 ;
        RECT 65.380 -118.120 65.720 -117.600 ;
        RECT 76.690 -118.300 76.990 -117.730 ;
      LAYER met2 ;
        RECT -63.710 -82.380 -62.120 -81.880 ;
        RECT -63.710 -84.340 40.000 -82.380 ;
        RECT -63.710 -232.700 -62.120 -84.340 ;
        RECT 37.250 -94.900 39.210 -84.340 ;
        RECT 35.450 -99.450 41.140 -94.900 ;
        RECT 65.080 -117.410 66.030 -116.840 ;
        RECT 76.260 -117.410 77.490 -117.120 ;
        RECT 65.080 -118.240 77.490 -117.410 ;
        RECT 65.080 -118.480 66.030 -118.240 ;
        RECT 76.260 -118.710 77.490 -118.240 ;
        RECT 28.480 -232.700 29.280 -232.550 ;
        RECT -63.710 -233.930 29.280 -232.700 ;
        RECT -63.360 -234.110 29.280 -233.930 ;
        RECT 28.480 -248.450 29.280 -234.110 ;
        RECT 41.580 -248.450 42.650 -248.360 ;
        RECT 28.480 -249.200 42.690 -248.450 ;
        RECT 41.580 -249.400 42.650 -249.200 ;
        RECT 41.420 -348.900 42.770 -249.400 ;
        RECT 41.840 -350.900 42.140 -348.900 ;
    END
  END AIN3
  PIN SEL2
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT 41.820 210.880 41.990 211.210 ;
        RECT 43.370 210.880 43.540 211.210 ;
        RECT 45.140 210.830 45.310 211.160 ;
        RECT 46.780 210.830 46.950 211.160 ;
        RECT 43.010 179.200 43.180 179.530 ;
        RECT 44.560 179.200 44.730 179.530 ;
        RECT 46.650 179.180 46.820 179.510 ;
        RECT 48.290 179.180 48.460 179.510 ;
      LAYER mcon ;
        RECT 41.820 210.960 41.990 211.130 ;
        RECT 43.370 210.960 43.540 211.130 ;
        RECT 45.140 210.910 45.310 211.080 ;
        RECT 46.780 210.910 46.950 211.080 ;
        RECT 43.010 179.280 43.180 179.450 ;
        RECT 44.560 179.280 44.730 179.450 ;
        RECT 46.650 179.260 46.820 179.430 ;
        RECT 48.290 179.260 48.460 179.430 ;
      LAYER met1 ;
        RECT 43.710 223.080 45.190 224.210 ;
        RECT 44.190 213.610 44.610 223.080 ;
        RECT 35.590 213.370 36.010 213.480 ;
        RECT 44.300 213.380 44.520 213.610 ;
        RECT 39.860 213.370 44.520 213.380 ;
        RECT 35.500 212.860 44.520 213.370 ;
        RECT 35.500 212.850 40.060 212.860 ;
        RECT 35.590 200.690 36.010 212.850 ;
        RECT 44.300 212.410 44.520 212.860 ;
        RECT 44.270 211.260 44.530 212.410 ;
        RECT 41.730 210.860 42.030 211.250 ;
        RECT 43.340 211.200 45.350 211.260 ;
        RECT 43.340 210.810 45.360 211.200 ;
        RECT 46.720 210.810 46.990 211.200 ;
        RECT 35.560 196.890 36.010 200.690 ;
        RECT 35.590 185.880 36.010 196.890 ;
        RECT 34.370 182.060 36.720 185.880 ;
        RECT 40.900 185.200 42.490 185.950 ;
        RECT 40.900 184.680 45.870 185.200 ;
        RECT 40.900 183.990 45.880 184.680 ;
        RECT 40.900 182.530 42.490 183.990 ;
        RECT 45.330 183.450 45.880 183.990 ;
        RECT 42.940 182.900 48.590 183.450 ;
        RECT 42.940 182.240 43.190 182.900 ;
        RECT 42.940 181.740 43.200 182.240 ;
        RECT 42.950 179.530 43.200 181.740 ;
        RECT 42.910 179.510 43.200 179.530 ;
        RECT 42.910 179.220 43.210 179.510 ;
        RECT 42.910 179.200 43.200 179.220 ;
        RECT 44.520 179.200 44.800 179.530 ;
        RECT 48.270 179.500 48.580 182.900 ;
        RECT 46.560 179.490 46.840 179.500 ;
        RECT 46.560 179.200 46.850 179.490 ;
        RECT 46.560 179.170 46.840 179.200 ;
        RECT 48.240 179.170 48.580 179.500 ;
        RECT 48.270 179.160 48.580 179.170 ;
      LAYER via ;
        RECT 44.190 223.480 44.490 223.760 ;
        RECT 35.030 183.540 35.700 184.840 ;
        RECT 41.440 184.070 41.830 185.030 ;
      LAYER met2 ;
        RECT 44.330 326.100 44.630 328.100 ;
        RECT 43.940 224.160 45.100 326.100 ;
        RECT 43.780 223.140 45.100 224.160 ;
        RECT 43.940 222.620 45.100 223.140 ;
        RECT 34.550 185.090 36.500 185.210 ;
        RECT 41.040 185.090 42.380 185.110 ;
        RECT 34.550 183.990 42.380 185.090 ;
        RECT 34.550 183.780 36.480 183.990 ;
        RECT 41.130 183.920 42.380 183.990 ;
        RECT 34.550 183.490 36.520 183.780 ;
        RECT 34.550 183.300 36.500 183.490 ;
    END
  END SEL2
  PIN DIGITALIN2
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT 42.740 196.030 42.910 196.360 ;
        RECT 44.290 196.030 44.460 196.360 ;
        RECT 46.510 196.050 46.680 196.380 ;
        RECT 48.150 196.050 48.320 196.380 ;
        RECT 42.900 175.740 43.070 176.070 ;
        RECT 44.450 175.740 44.620 176.070 ;
        RECT 46.670 175.760 46.840 176.090 ;
        RECT 48.310 175.760 48.480 176.090 ;
      LAYER mcon ;
        RECT 42.740 196.110 42.910 196.280 ;
        RECT 44.290 196.110 44.460 196.280 ;
        RECT 46.510 196.130 46.680 196.300 ;
        RECT 48.150 196.130 48.320 196.300 ;
        RECT 42.900 175.820 43.070 175.990 ;
        RECT 44.450 175.820 44.620 175.990 ;
        RECT 46.670 175.840 46.840 176.010 ;
        RECT 48.310 175.840 48.480 176.010 ;
      LAYER met1 ;
        RECT 42.670 196.030 42.950 196.360 ;
        RECT 44.250 194.130 44.530 196.370 ;
        RECT 46.430 196.050 46.710 196.380 ;
        RECT 44.230 194.070 44.530 194.130 ;
        RECT 48.120 194.070 48.470 196.410 ;
        RECT 51.160 194.620 52.380 194.660 ;
        RECT 44.230 194.040 48.920 194.070 ;
        RECT 49.290 194.040 49.870 194.350 ;
        RECT 44.230 193.590 49.870 194.040 ;
        RECT 44.230 193.570 48.920 193.590 ;
        RECT 44.230 193.530 44.520 193.570 ;
        RECT 49.290 193.390 49.870 193.590 ;
        RECT 50.960 193.380 52.380 194.620 ;
        RECT 51.160 191.670 52.380 193.380 ;
        RECT 61.160 184.680 63.860 184.970 ;
        RECT 59.790 181.890 63.860 184.680 ;
        RECT 61.160 181.610 63.860 181.890 ;
        RECT 42.830 175.740 43.110 176.070 ;
        RECT 44.410 173.840 44.690 176.080 ;
        RECT 46.590 175.760 46.870 176.090 ;
        RECT 44.390 173.780 44.690 173.840 ;
        RECT 48.280 173.780 48.630 176.120 ;
        RECT 51.250 174.330 52.590 174.620 ;
        RECT 44.390 173.750 49.080 173.780 ;
        RECT 49.450 173.750 50.030 174.060 ;
        RECT 44.390 173.300 50.030 173.750 ;
        RECT 44.390 173.280 49.080 173.300 ;
        RECT 44.390 173.240 44.680 173.280 ;
        RECT 49.450 173.100 50.030 173.300 ;
        RECT 51.120 173.090 52.590 174.330 ;
        RECT 51.250 172.130 52.590 173.090 ;
      LAYER via ;
        RECT 49.460 193.700 49.720 194.130 ;
        RECT 51.230 193.850 51.490 194.290 ;
        RECT 51.560 192.590 51.950 194.190 ;
        RECT 60.270 182.570 60.830 184.280 ;
        RECT 62.280 182.740 62.940 183.760 ;
        RECT 49.620 173.410 49.880 173.840 ;
        RECT 51.390 173.560 51.650 174.000 ;
        RECT 51.760 173.060 52.020 174.100 ;
      LAYER met2 ;
        RECT 47.090 326.100 47.390 328.090 ;
        RECT 46.920 222.770 47.590 326.100 ;
        RECT 45.880 222.310 47.610 222.770 ;
        RECT 45.900 219.100 46.520 222.310 ;
        RECT 46.920 222.300 47.590 222.310 ;
        RECT 45.900 218.250 63.170 219.100 ;
        RECT 62.160 196.500 63.050 218.250 ;
        RECT 62.110 196.380 63.050 196.500 ;
        RECT 51.050 194.510 51.680 194.530 ;
        RECT 49.370 194.200 49.790 194.260 ;
        RECT 51.050 194.250 52.270 194.510 ;
        RECT 53.880 194.250 54.140 194.370 ;
        RECT 51.050 194.200 54.140 194.250 ;
        RECT 49.370 193.630 54.140 194.200 ;
        RECT 49.370 193.490 49.790 193.630 ;
        RECT 51.050 193.460 54.140 193.630 ;
        RECT 51.360 192.460 54.140 193.460 ;
        RECT 51.360 191.850 52.270 192.460 ;
        RECT 53.880 184.020 54.140 192.460 ;
        RECT 62.110 184.710 63.000 196.380 ;
        RECT 59.970 184.020 61.210 184.510 ;
        RECT 53.880 183.210 61.210 184.020 ;
        RECT 53.880 182.310 54.160 183.210 ;
        RECT 59.980 182.530 61.210 183.210 ;
        RECT 51.420 174.240 52.360 174.460 ;
        RECT 51.210 174.060 52.360 174.240 ;
        RECT 53.880 174.060 54.140 182.310 ;
        RECT 60.010 182.050 61.210 182.530 ;
        RECT 61.620 181.770 63.700 184.710 ;
        RECT 49.530 173.910 49.950 173.970 ;
        RECT 51.210 173.910 54.140 174.060 ;
        RECT 49.530 173.370 54.140 173.910 ;
        RECT 49.530 173.340 54.120 173.370 ;
        RECT 49.530 173.200 49.950 173.340 ;
        RECT 51.210 173.170 54.120 173.340 ;
        RECT 51.420 172.790 54.120 173.170 ;
        RECT 51.420 172.440 52.360 172.790 ;
    END
  END DIGITALIN2
  PIN AIN2
    ANTENNADIFFAREA 23.199999 ;
    PORT
      LAYER li1 ;
        RECT 65.425 87.780 85.465 87.950 ;
        RECT -1.135 86.490 18.905 86.660 ;
        RECT 65.230 83.340 85.270 83.510 ;
        RECT -1.330 82.050 18.710 82.220 ;
      LAYER mcon ;
        RECT 65.505 87.780 85.385 87.950 ;
        RECT -1.055 86.490 18.825 86.660 ;
        RECT 65.310 83.340 85.190 83.510 ;
        RECT -1.250 82.050 18.630 82.220 ;
      LAYER met1 ;
        RECT 62.550 91.920 63.740 92.670 ;
        RECT 18.140 91.850 63.740 91.920 ;
        RECT 18.090 91.570 63.740 91.850 ;
        RECT 18.090 89.340 18.490 91.570 ;
        RECT 17.940 88.960 18.850 89.340 ;
        RECT 17.940 88.940 21.880 88.960 ;
        RECT 17.940 88.570 21.890 88.940 ;
        RECT 17.930 88.250 21.890 88.570 ;
        RECT 17.930 87.230 18.850 88.250 ;
        RECT 17.930 86.690 18.840 87.230 ;
        RECT -1.115 86.460 18.885 86.690 ;
        RECT -1.310 82.020 18.690 82.250 ;
        RECT 18.250 80.960 18.600 82.020 ;
        RECT 21.200 80.960 21.890 88.250 ;
        RECT 18.140 80.110 21.890 80.960 ;
        RECT 18.140 80.100 21.770 80.110 ;
        RECT 35.110 74.170 36.500 91.570 ;
        RECT 62.550 90.760 63.740 91.570 ;
        RECT 73.770 92.620 75.130 92.890 ;
        RECT 85.060 92.620 85.410 92.690 ;
        RECT 73.770 91.740 85.410 92.620 ;
        RECT 73.770 91.090 75.130 91.740 ;
        RECT 85.060 90.630 85.410 91.740 ;
        RECT 84.500 90.250 85.410 90.630 ;
        RECT 84.500 90.230 88.440 90.250 ;
        RECT 84.500 89.860 88.450 90.230 ;
        RECT 84.490 89.540 88.450 89.860 ;
        RECT 84.490 88.520 85.410 89.540 ;
        RECT 84.490 87.980 85.400 88.520 ;
        RECT 65.445 87.750 85.445 87.980 ;
        RECT 65.250 83.310 85.250 83.540 ;
        RECT 84.810 82.250 85.160 83.310 ;
        RECT 87.760 82.250 88.450 89.540 ;
        RECT 84.700 81.400 88.450 82.250 ;
        RECT 84.700 81.390 88.330 81.400 ;
        RECT 32.330 68.400 39.510 74.170 ;
      LAYER via ;
        RECT 62.960 91.710 63.300 92.230 ;
        RECT 74.270 91.840 74.570 92.410 ;
        RECT 35.260 70.470 36.580 72.390 ;
      LAYER met2 ;
        RECT 39.740 326.100 40.040 328.100 ;
        RECT 39.290 224.560 40.440 326.100 ;
        RECT 39.160 223.930 40.440 224.560 ;
        RECT 39.160 223.310 40.230 223.930 ;
        RECT 26.060 222.560 40.270 223.310 ;
        RECT 26.060 208.220 26.860 222.560 ;
        RECT 39.160 222.470 40.230 222.560 ;
        RECT -65.780 208.040 26.860 208.220 ;
        RECT -66.130 206.810 26.860 208.040 ;
        RECT -66.130 58.450 -64.540 206.810 ;
        RECT 26.060 206.660 26.860 206.810 ;
        RECT 62.660 92.350 63.610 92.590 ;
        RECT 73.840 92.350 75.070 92.820 ;
        RECT 62.660 91.520 75.070 92.350 ;
        RECT 62.660 90.950 63.610 91.520 ;
        RECT 73.840 91.230 75.070 91.520 ;
        RECT 33.030 69.010 38.720 73.560 ;
        RECT 34.830 58.450 36.790 69.010 ;
        RECT -66.130 56.490 37.580 58.450 ;
        RECT -66.130 55.990 -64.540 56.490 ;
    END
  END AIN2
  PIN vssa1
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT -315.150 -273.900 -305.150 251.100 ;
        RECT 154.850 -273.900 164.850 251.100 ;
      LAYER via2 ;
        RECT -312.650 243.600 -307.650 248.600 ;
        RECT -312.650 -271.400 -307.650 -266.400 ;
        RECT 157.350 243.600 162.350 248.600 ;
        RECT 157.350 -271.400 162.350 -266.400 ;
      LAYER met3 ;
        RECT -400.150 241.100 249.850 251.100 ;
        RECT -400.150 -273.900 249.850 -263.900 ;
    END
  END vssa1
  PIN vdda1
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 15.150 135.040 38.120 138.120 ;
        RECT 93.080 134.610 116.050 137.690 ;
        RECT 15.210 128.850 38.180 131.930 ;
        RECT 93.140 128.420 116.110 131.500 ;
        RECT -2.600 84.640 20.370 87.720 ;
        RECT 63.960 85.930 86.930 89.010 ;
        RECT 0.990 35.840 23.960 38.920 ;
        RECT 65.810 38.830 88.780 41.910 ;
        RECT -214.290 -11.280 -211.210 11.690 ;
        RECT -208.100 -11.340 -205.020 11.630 ;
        RECT -163.890 6.470 -160.810 29.440 ;
        RECT -115.090 2.880 -112.010 25.850 ;
        RECT -165.180 -60.090 -162.100 -37.120 ;
        RECT -118.080 -61.940 -115.000 -38.970 ;
        RECT 3.410 -64.810 26.380 -61.730 ;
        RECT -213.860 -89.210 -210.780 -66.240 ;
        RECT -207.670 -89.270 -204.590 -66.300 ;
        RECT 68.230 -67.800 91.200 -64.720 ;
        RECT -0.180 -113.610 22.790 -110.530 ;
        RECT 66.380 -114.900 89.350 -111.820 ;
        RECT 17.630 -157.820 40.600 -154.740 ;
        RECT 95.560 -157.390 118.530 -154.310 ;
        RECT 17.570 -164.010 40.540 -160.930 ;
        RECT 95.500 -163.580 118.470 -160.500 ;
      LAYER li1 ;
        RECT -11.400 143.030 8.640 143.200 ;
        RECT 66.530 142.600 86.570 142.770 ;
        RECT 15.540 137.560 37.730 137.730 ;
        RECT 15.540 135.600 15.710 137.560 ;
        RECT 16.615 136.100 36.655 136.270 ;
        RECT 37.560 135.600 37.730 137.560 ;
        RECT 15.540 135.430 37.730 135.600 ;
        RECT 93.470 137.130 115.660 137.300 ;
        RECT 35.750 135.420 36.550 135.430 ;
        RECT 93.470 135.170 93.640 137.130 ;
        RECT 94.545 135.670 114.585 135.840 ;
        RECT 115.490 135.170 115.660 137.130 ;
        RECT 93.470 135.000 115.660 135.170 ;
        RECT 113.680 134.990 114.480 135.000 ;
        RECT 35.800 131.540 36.520 131.550 ;
        RECT 15.600 131.370 37.790 131.540 ;
        RECT 15.600 129.410 15.770 131.370 ;
        RECT 35.800 131.350 36.520 131.370 ;
        RECT 16.675 130.700 36.715 130.870 ;
        RECT 37.620 129.410 37.790 131.370 ;
        RECT 113.730 131.110 114.450 131.120 ;
        RECT 15.600 129.240 37.790 129.410 ;
        RECT 93.530 130.940 115.720 131.110 ;
        RECT 93.530 128.980 93.700 130.940 ;
        RECT 113.730 130.920 114.450 130.940 ;
        RECT 94.605 130.270 114.645 130.440 ;
        RECT 115.550 128.980 115.720 130.940 ;
        RECT 93.530 128.810 115.720 128.980 ;
        RECT -11.660 124.250 8.380 124.420 ;
        RECT 66.270 123.820 86.310 123.990 ;
        RECT 64.350 88.450 86.540 88.620 ;
        RECT -2.210 87.160 19.980 87.330 ;
        RECT -2.210 85.200 -2.040 87.160 ;
        RECT 19.810 85.200 19.980 87.160 ;
        RECT 64.350 86.490 64.520 88.450 ;
        RECT 86.370 86.490 86.540 88.450 ;
        RECT 64.350 86.320 86.540 86.490 ;
        RECT -2.210 85.030 19.980 85.200 ;
        RECT 66.200 41.350 88.390 41.520 ;
        RECT 66.200 39.390 66.370 41.350 ;
        RECT 88.220 39.390 88.390 41.350 ;
        RECT 66.200 39.220 88.390 39.390 ;
        RECT -219.370 18.200 -219.200 38.240 ;
        RECT -200.590 18.460 -200.420 38.500 ;
        RECT 1.380 38.360 23.570 38.530 ;
        RECT 1.380 36.400 1.550 38.360 ;
        RECT 23.400 36.400 23.570 38.360 ;
        RECT 1.380 36.230 23.570 36.400 ;
        RECT -163.500 28.880 -161.200 29.050 ;
        RECT -213.900 11.130 -211.600 11.300 ;
        RECT -213.900 -10.720 -213.730 11.130 ;
        RECT -212.440 -9.815 -212.270 10.225 ;
        RECT -211.770 -8.910 -211.600 11.130 ;
        RECT -207.710 11.070 -205.410 11.240 ;
        RECT -211.770 -9.710 -211.590 -8.910 ;
        RECT -207.710 -8.960 -207.540 11.070 ;
        RECT -207.720 -9.680 -207.520 -8.960 ;
        RECT -211.770 -10.720 -211.600 -9.710 ;
        RECT -213.900 -10.890 -211.600 -10.720 ;
        RECT -207.710 -10.780 -207.540 -9.680 ;
        RECT -207.040 -9.875 -206.870 10.165 ;
        RECT -205.580 -10.780 -205.410 11.070 ;
        RECT -163.500 7.030 -163.330 28.880 ;
        RECT -161.370 7.030 -161.200 28.880 ;
        RECT -163.500 6.860 -161.200 7.030 ;
        RECT -114.700 25.290 -112.400 25.460 ;
        RECT -114.700 3.440 -114.530 25.290 ;
        RECT -112.570 3.440 -112.400 25.290 ;
        RECT -114.700 3.270 -112.400 3.440 ;
        RECT -207.710 -10.950 -205.410 -10.780 ;
        RECT -164.790 -37.680 -162.490 -37.510 ;
        RECT -218.940 -59.730 -218.770 -39.690 ;
        RECT -200.160 -59.470 -199.990 -39.430 ;
        RECT -164.790 -59.530 -164.620 -37.680 ;
        RECT -162.660 -59.530 -162.490 -37.680 ;
        RECT -164.790 -59.700 -162.490 -59.530 ;
        RECT -117.690 -39.530 -115.390 -39.360 ;
        RECT -117.690 -61.380 -117.520 -39.530 ;
        RECT -115.560 -61.380 -115.390 -39.530 ;
        RECT -117.690 -61.550 -115.390 -61.380 ;
        RECT 3.800 -62.290 25.990 -62.120 ;
        RECT 3.800 -64.250 3.970 -62.290 ;
        RECT 25.820 -64.250 25.990 -62.290 ;
        RECT 3.800 -64.420 25.990 -64.250 ;
        RECT 68.620 -65.280 90.810 -65.110 ;
        RECT -213.470 -66.800 -211.170 -66.630 ;
        RECT -213.470 -88.650 -213.300 -66.800 ;
        RECT -212.010 -87.745 -211.840 -67.705 ;
        RECT -211.340 -86.840 -211.170 -66.800 ;
        RECT -207.280 -66.860 -204.980 -66.690 ;
        RECT -211.340 -87.640 -211.160 -86.840 ;
        RECT -207.280 -86.890 -207.110 -66.860 ;
        RECT -207.290 -87.610 -207.090 -86.890 ;
        RECT -211.340 -88.650 -211.170 -87.640 ;
        RECT -213.470 -88.820 -211.170 -88.650 ;
        RECT -207.280 -88.710 -207.110 -87.610 ;
        RECT -206.610 -87.805 -206.440 -67.765 ;
        RECT -205.150 -88.710 -204.980 -66.860 ;
        RECT 68.620 -67.240 68.790 -65.280 ;
        RECT 90.640 -67.240 90.810 -65.280 ;
        RECT 68.620 -67.410 90.810 -67.240 ;
        RECT -207.280 -88.880 -204.980 -88.710 ;
        RECT 0.210 -111.090 22.400 -110.920 ;
        RECT 0.210 -113.050 0.380 -111.090 ;
        RECT 22.230 -113.050 22.400 -111.090 ;
        RECT 0.210 -113.220 22.400 -113.050 ;
        RECT 66.770 -112.380 88.960 -112.210 ;
        RECT 66.770 -114.340 66.940 -112.380 ;
        RECT 88.790 -114.340 88.960 -112.380 ;
        RECT 66.770 -114.510 88.960 -114.340 ;
        RECT 68.690 -149.880 88.730 -149.710 ;
        RECT -9.240 -150.310 10.800 -150.140 ;
        RECT 95.950 -154.870 118.140 -154.700 ;
        RECT 18.020 -155.300 40.210 -155.130 ;
        RECT 18.020 -157.260 18.190 -155.300 ;
        RECT 19.095 -156.760 39.135 -156.590 ;
        RECT 38.220 -157.260 38.940 -157.240 ;
        RECT 40.040 -157.260 40.210 -155.300 ;
        RECT 95.950 -156.830 96.120 -154.870 ;
        RECT 97.025 -156.330 117.065 -156.160 ;
        RECT 116.150 -156.830 116.870 -156.810 ;
        RECT 117.970 -156.830 118.140 -154.870 ;
        RECT 95.950 -157.000 118.140 -156.830 ;
        RECT 116.150 -157.010 116.870 -157.000 ;
        RECT 18.020 -157.430 40.210 -157.260 ;
        RECT 38.220 -157.440 38.940 -157.430 ;
        RECT 116.100 -160.890 116.900 -160.880 ;
        RECT 95.890 -161.060 118.080 -160.890 ;
        RECT 38.170 -161.320 38.970 -161.310 ;
        RECT 17.960 -161.490 40.150 -161.320 ;
        RECT 17.960 -163.450 18.130 -161.490 ;
        RECT 19.035 -162.160 39.075 -161.990 ;
        RECT 39.980 -163.450 40.150 -161.490 ;
        RECT 95.890 -163.020 96.060 -161.060 ;
        RECT 96.965 -161.730 117.005 -161.560 ;
        RECT 117.910 -163.020 118.080 -161.060 ;
        RECT 95.890 -163.190 118.080 -163.020 ;
        RECT 17.960 -163.620 40.150 -163.450 ;
        RECT 68.950 -168.660 88.990 -168.490 ;
        RECT -8.980 -169.090 11.060 -168.920 ;
      LAYER mcon ;
        RECT -11.320 143.030 8.560 143.200 ;
        RECT 66.610 142.600 86.490 142.770 ;
        RECT 16.695 136.100 36.575 136.270 ;
        RECT 94.625 135.670 114.505 135.840 ;
        RECT 16.755 130.700 36.635 130.870 ;
        RECT 94.685 130.270 114.565 130.440 ;
        RECT -11.580 124.250 8.300 124.420 ;
        RECT 66.350 123.820 86.230 123.990 ;
        RECT 65.370 88.450 65.970 88.620 ;
        RECT -1.190 87.160 -0.590 87.330 ;
        RECT 67.220 41.350 67.820 41.520 ;
        RECT -219.370 18.280 -219.200 38.160 ;
        RECT -200.590 18.540 -200.420 38.420 ;
        RECT 2.400 38.360 3.000 38.530 ;
        RECT -163.500 27.430 -163.330 28.030 ;
        RECT -212.440 -9.735 -212.270 10.145 ;
        RECT -211.770 -9.710 -211.590 -8.910 ;
        RECT -207.720 -9.680 -207.520 -8.960 ;
        RECT -207.040 -9.795 -206.870 10.085 ;
        RECT -114.700 23.840 -114.530 24.440 ;
        RECT -164.790 -39.130 -164.620 -38.530 ;
        RECT -218.940 -59.650 -218.770 -39.770 ;
        RECT -200.160 -59.390 -199.990 -39.510 ;
        RECT -117.690 -40.980 -117.520 -40.380 ;
        RECT 4.820 -64.420 5.420 -64.250 ;
        RECT -212.010 -87.665 -211.840 -67.785 ;
        RECT -211.340 -87.640 -211.160 -86.840 ;
        RECT -207.290 -87.610 -207.090 -86.890 ;
        RECT -206.610 -87.725 -206.440 -67.845 ;
        RECT 69.640 -67.410 70.240 -67.240 ;
        RECT 1.230 -113.220 1.830 -113.050 ;
        RECT 67.790 -114.510 68.390 -114.340 ;
        RECT 68.770 -149.880 88.650 -149.710 ;
        RECT -9.160 -150.310 10.720 -150.140 ;
        RECT 19.175 -156.760 39.055 -156.590 ;
        RECT 97.105 -156.330 116.985 -156.160 ;
        RECT 116.100 -161.060 116.900 -160.880 ;
        RECT 38.170 -161.490 38.970 -161.310 ;
        RECT 19.115 -162.160 38.995 -161.990 ;
        RECT 97.045 -161.730 116.925 -161.560 ;
        RECT 69.030 -168.660 88.910 -168.490 ;
        RECT -8.900 -169.090 10.980 -168.920 ;
      LAYER met1 ;
        RECT 10.610 146.060 10.990 146.070 ;
        RECT 48.150 146.060 48.640 146.080 ;
        RECT 8.260 145.390 48.640 146.060 ;
        RECT 88.540 145.630 88.920 145.640 ;
        RECT 126.080 145.630 126.570 145.650 ;
        RECT 8.260 143.230 8.570 145.390 ;
        RECT -11.380 143.000 8.620 143.230 ;
        RECT 16.635 136.070 36.635 136.300 ;
        RECT 35.730 135.660 36.560 136.070 ;
        RECT 35.560 135.360 36.620 135.660 ;
        RECT 35.730 134.330 36.560 135.360 ;
        RECT 48.150 135.160 48.640 145.390 ;
        RECT 86.190 144.960 126.570 145.630 ;
        RECT 86.190 142.800 86.500 144.960 ;
        RECT 66.550 142.570 86.550 142.800 ;
        RECT 94.565 135.640 114.565 135.870 ;
        RECT 113.660 135.230 114.490 135.640 ;
        RECT 50.550 135.160 51.240 135.180 ;
        RECT 48.150 134.330 51.240 135.160 ;
        RECT 113.490 134.930 114.550 135.230 ;
        RECT 35.730 134.060 51.240 134.330 ;
        RECT 35.730 132.250 48.640 134.060 ;
        RECT 35.730 130.900 36.560 132.250 ;
        RECT 16.695 130.670 36.695 130.900 ;
        RECT -11.640 124.220 8.360 124.450 ;
        RECT 7.690 124.040 8.310 124.220 ;
        RECT 7.690 123.250 8.320 124.040 ;
        RECT 7.700 119.160 8.250 123.250 ;
        RECT 48.150 119.160 48.640 132.250 ;
        RECT 7.660 118.140 48.690 119.160 ;
        RECT 48.150 118.110 48.640 118.140 ;
        RECT 50.550 115.610 51.240 134.060 ;
        RECT 113.660 133.900 114.490 134.930 ;
        RECT 126.080 134.580 126.570 144.960 ;
        RECT 126.790 134.580 141.240 134.710 ;
        RECT 126.080 133.950 141.240 134.580 ;
        RECT 126.080 133.900 127.260 133.950 ;
        RECT 113.660 133.880 127.260 133.900 ;
        RECT 113.660 131.820 126.570 133.880 ;
        RECT 113.660 130.470 114.490 131.820 ;
        RECT 94.625 130.240 114.625 130.470 ;
        RECT 66.290 123.790 86.290 124.020 ;
        RECT 85.620 123.610 86.240 123.790 ;
        RECT 85.620 122.820 86.250 123.610 ;
        RECT 85.630 118.730 86.180 122.820 ;
        RECT 126.080 118.730 126.570 131.820 ;
        RECT 140.730 123.960 141.240 133.950 ;
        RECT 140.710 122.700 141.270 123.960 ;
        RECT 85.590 117.710 126.620 118.730 ;
        RECT 140.730 118.330 141.240 122.700 ;
        RECT 148.160 118.340 150.390 118.400 ;
        RECT 147.230 118.330 150.390 118.340 ;
        RECT 126.080 117.680 126.570 117.710 ;
        RECT 50.530 114.890 51.240 115.610 ;
        RECT 140.730 117.470 150.390 118.330 ;
        RECT 50.530 97.230 51.220 114.890 ;
        RECT -1.410 96.910 51.450 97.230 ;
        RECT 140.730 97.030 141.240 117.470 ;
        RECT 138.640 96.910 141.240 97.030 ;
        RECT -1.410 96.250 141.240 96.910 ;
        RECT -1.290 87.960 -0.550 96.250 ;
        RECT 50.390 95.310 141.240 96.250 ;
        RECT 50.390 95.290 140.730 95.310 ;
        RECT 50.390 95.230 139.110 95.290 ;
        RECT 65.380 89.470 65.940 95.230 ;
        RECT 65.360 88.690 66.010 89.470 ;
        RECT 65.300 88.390 66.020 88.690 ;
        RECT -1.200 87.400 -0.550 87.960 ;
        RECT -1.260 87.100 -0.540 87.400 ;
        RECT 104.190 54.490 105.490 95.230 ;
        RECT 67.100 53.900 105.650 54.490 ;
        RECT 67.110 52.350 67.890 53.900 ;
        RECT 2.260 50.910 67.890 52.350 ;
        RECT 2.350 38.890 3.130 50.910 ;
        RECT 67.110 41.850 67.890 50.910 ;
        RECT 67.210 41.590 67.860 41.850 ;
        RECT 67.150 41.290 67.870 41.590 ;
        RECT 2.390 38.600 3.040 38.890 ;
        RECT -219.400 18.580 -219.170 38.220 ;
        RECT -222.230 18.270 -219.170 18.580 ;
        RECT -200.620 19.150 -200.390 38.480 ;
        RECT 2.330 38.300 3.050 38.600 ;
        RECT -173.400 28.130 -172.420 28.250 ;
        RECT -173.400 28.040 -164.130 28.130 ;
        RECT -163.570 28.040 -163.270 28.100 ;
        RECT -173.400 27.390 -163.270 28.040 ;
        RECT -200.620 19.140 -199.420 19.150 ;
        RECT -195.330 19.140 -194.310 19.180 ;
        RECT -200.620 18.590 -194.310 19.140 ;
        RECT -200.620 18.530 -199.420 18.590 ;
        RECT -200.620 18.480 -200.390 18.530 ;
        RECT -200.210 18.520 -199.420 18.530 ;
        RECT -222.230 16.230 -221.560 18.270 ;
        RECT -219.400 18.220 -219.170 18.270 ;
        RECT -222.240 15.850 -221.560 16.230 ;
        RECT -222.230 -21.310 -221.560 15.850 ;
        RECT -212.470 -8.890 -212.240 10.205 ;
        RECT -211.830 -8.890 -211.530 -8.720 ;
        RECT -207.070 -8.890 -206.840 10.145 ;
        RECT -212.470 -9.720 -206.840 -8.890 ;
        RECT -212.470 -9.795 -212.240 -9.720 ;
        RECT -211.830 -9.780 -211.530 -9.720 ;
        RECT -210.500 -21.310 -208.420 -9.720 ;
        RECT -207.070 -9.855 -206.840 -9.720 ;
        RECT -195.330 -21.310 -194.310 18.590 ;
        RECT -222.250 -21.800 -194.280 -21.310 ;
        RECT -211.330 -23.710 -210.230 -21.800 ;
        RECT -195.330 -21.850 -194.310 -21.800 ;
        RECT -173.400 -23.550 -172.420 27.390 ;
        RECT -163.570 27.380 -163.270 27.390 ;
        RECT -128.520 24.490 -127.080 24.580 ;
        RECT -128.520 24.450 -115.060 24.490 ;
        RECT -114.770 24.450 -114.470 24.510 ;
        RECT -128.520 23.800 -114.470 24.450 ;
        RECT -128.520 23.710 -115.060 23.800 ;
        RECT -114.770 23.790 -114.470 23.800 ;
        RECT -173.400 -23.690 -171.400 -23.550 ;
        RECT -191.780 -23.710 -171.400 -23.690 ;
        RECT -211.350 -24.380 -171.400 -23.710 ;
        RECT -211.350 -24.400 -191.060 -24.380 ;
        RECT -173.400 -24.610 -171.400 -24.380 ;
        RECT -173.080 -38.540 -171.400 -24.610 ;
        RECT -164.860 -38.520 -164.560 -38.460 ;
        RECT -165.640 -38.540 -164.560 -38.520 ;
        RECT -173.080 -39.100 -164.560 -38.540 ;
        RECT -218.970 -59.350 -218.740 -39.710 ;
        RECT -221.800 -59.660 -218.740 -59.350 ;
        RECT -200.190 -58.780 -199.960 -39.450 ;
        RECT -200.190 -58.790 -198.990 -58.780 ;
        RECT -194.900 -58.790 -193.880 -58.750 ;
        RECT -200.190 -59.340 -193.880 -58.790 ;
        RECT -200.190 -59.400 -198.990 -59.340 ;
        RECT -200.190 -59.450 -199.960 -59.400 ;
        RECT -199.780 -59.410 -198.990 -59.400 ;
        RECT -221.800 -61.700 -221.130 -59.660 ;
        RECT -218.970 -59.710 -218.740 -59.660 ;
        RECT -221.810 -62.080 -221.130 -61.700 ;
        RECT -221.800 -99.240 -221.130 -62.080 ;
        RECT -212.040 -86.820 -211.810 -67.725 ;
        RECT -211.400 -86.820 -211.100 -86.650 ;
        RECT -206.640 -86.820 -206.410 -67.785 ;
        RECT -212.040 -87.650 -206.410 -86.820 ;
        RECT -212.040 -87.725 -211.810 -87.650 ;
        RECT -211.400 -87.710 -211.100 -87.650 ;
        RECT -210.070 -99.240 -207.990 -87.650 ;
        RECT -206.640 -87.785 -206.410 -87.650 ;
        RECT -194.900 -99.240 -193.880 -59.340 ;
        RECT -173.080 -77.350 -171.400 -39.100 ;
        RECT -165.640 -39.170 -164.560 -39.100 ;
        RECT -164.860 -39.180 -164.560 -39.170 ;
        RECT -130.660 -40.270 -130.070 -40.260 ;
        RECT -128.520 -40.270 -127.080 23.710 ;
        RECT -130.660 -40.370 -118.020 -40.270 ;
        RECT -117.760 -40.370 -117.460 -40.310 ;
        RECT -130.660 -41.020 -117.460 -40.370 ;
        RECT -130.660 -41.050 -118.020 -41.020 ;
        RECT -117.760 -41.030 -117.460 -41.020 ;
        RECT -130.660 -77.350 -130.070 -41.050 ;
        RECT 4.750 -64.490 5.470 -64.190 ;
        RECT 4.810 -64.780 5.460 -64.490 ;
        RECT 4.770 -76.800 5.550 -64.780 ;
        RECT 69.570 -67.480 70.290 -67.180 ;
        RECT 69.630 -67.740 70.280 -67.480 ;
        RECT 69.530 -76.800 70.310 -67.740 ;
        RECT -173.080 -78.650 -130.070 -77.350 ;
        RECT 4.680 -78.240 70.310 -76.800 ;
        RECT -221.820 -99.730 -193.850 -99.240 ;
        RECT -210.750 -99.950 -210.050 -99.730 ;
        RECT -194.900 -99.780 -193.880 -99.730 ;
        RECT -210.880 -100.420 -210.050 -99.950 ;
        RECT -210.880 -113.890 -210.120 -100.420 ;
        RECT -173.080 -111.800 -171.400 -78.650 ;
        RECT -130.660 -78.810 -130.070 -78.650 ;
        RECT 69.530 -79.790 70.310 -78.240 ;
        RECT 69.520 -80.380 108.070 -79.790 ;
        RECT -173.200 -112.270 -171.400 -111.800 ;
        RECT -200.130 -113.890 -198.870 -113.870 ;
        RECT -173.200 -113.890 -171.460 -112.270 ;
        RECT 1.160 -113.290 1.880 -112.990 ;
        RECT 1.220 -113.850 1.870 -113.290 ;
        RECT -210.880 -114.400 -171.480 -113.890 ;
        RECT -200.130 -114.430 -198.870 -114.400 ;
        RECT -194.500 -119.940 -193.640 -114.400 ;
        RECT -195.220 -121.540 -193.200 -119.940 ;
        RECT 1.130 -122.140 1.870 -113.850 ;
        RECT 67.720 -114.580 68.440 -114.280 ;
        RECT 67.780 -115.360 68.430 -114.580 ;
        RECT 67.800 -121.120 68.360 -115.360 ;
        RECT 106.610 -121.120 107.910 -80.380 ;
        RECT 52.810 -121.180 141.530 -121.120 ;
        RECT 52.810 -121.200 143.150 -121.180 ;
        RECT 52.810 -122.140 143.660 -121.200 ;
        RECT 1.010 -122.800 143.660 -122.140 ;
        RECT 1.010 -123.120 53.870 -122.800 ;
        RECT 141.060 -122.920 143.660 -122.800 ;
        RECT 52.950 -140.780 53.640 -123.120 ;
        RECT 52.950 -141.500 53.660 -140.780 ;
        RECT 50.570 -144.030 51.060 -144.000 ;
        RECT 10.080 -145.050 51.110 -144.030 ;
        RECT 10.120 -149.140 10.670 -145.050 ;
        RECT 10.110 -149.930 10.740 -149.140 ;
        RECT 10.110 -150.110 10.730 -149.930 ;
        RECT -9.220 -150.340 10.780 -150.110 ;
        RECT 19.115 -156.790 39.115 -156.560 ;
        RECT 38.150 -158.140 38.980 -156.790 ;
        RECT 50.570 -158.140 51.060 -145.050 ;
        RECT 38.150 -159.950 51.060 -158.140 ;
        RECT 52.970 -159.950 53.660 -141.500 ;
        RECT 143.150 -143.360 143.660 -122.920 ;
        RECT 148.160 -142.330 150.390 117.470 ;
        RECT 148.140 -143.360 150.450 -142.330 ;
        RECT 128.500 -143.600 128.990 -143.570 ;
        RECT 88.010 -144.620 129.040 -143.600 ;
        RECT 143.150 -144.220 150.450 -143.360 ;
        RECT 88.050 -148.710 88.600 -144.620 ;
        RECT 88.040 -149.500 88.670 -148.710 ;
        RECT 88.040 -149.680 88.660 -149.500 ;
        RECT 68.710 -149.910 88.710 -149.680 ;
        RECT 97.045 -156.360 117.045 -156.130 ;
        RECT 38.150 -160.220 53.660 -159.950 ;
        RECT 38.150 -161.250 38.980 -160.220 ;
        RECT 50.570 -161.050 53.660 -160.220 ;
        RECT 116.080 -157.710 116.910 -156.360 ;
        RECT 128.500 -157.710 128.990 -144.620 ;
        RECT 143.150 -148.590 143.660 -144.220 ;
        RECT 143.130 -149.850 143.690 -148.590 ;
        RECT 116.080 -159.770 128.990 -157.710 ;
        RECT 116.080 -159.790 129.680 -159.770 ;
        RECT 116.080 -160.820 116.910 -159.790 ;
        RECT 128.500 -159.840 129.680 -159.790 ;
        RECT 143.150 -159.840 143.660 -149.850 ;
        RECT 128.500 -160.470 143.660 -159.840 ;
        RECT 37.980 -161.550 39.040 -161.250 ;
        RECT 38.150 -161.960 38.980 -161.550 ;
        RECT 19.055 -162.190 39.055 -161.960 ;
        RECT -8.960 -169.120 11.040 -168.890 ;
        RECT 10.680 -171.280 10.990 -169.120 ;
        RECT 50.570 -171.280 51.060 -161.050 ;
        RECT 52.970 -161.070 53.660 -161.050 ;
        RECT 115.910 -161.120 116.970 -160.820 ;
        RECT 116.080 -161.530 116.910 -161.120 ;
        RECT 96.985 -161.760 116.985 -161.530 ;
        RECT 68.970 -168.690 88.970 -168.460 ;
        RECT 10.680 -171.950 51.060 -171.280 ;
        RECT 88.610 -170.850 88.920 -168.690 ;
        RECT 128.500 -170.850 128.990 -160.470 ;
        RECT 129.210 -160.600 143.660 -160.470 ;
        RECT 88.610 -171.520 128.990 -170.850 ;
        RECT 90.960 -171.530 91.340 -171.520 ;
        RECT 128.500 -171.540 128.990 -171.520 ;
        RECT 13.030 -171.960 13.410 -171.950 ;
        RECT 50.570 -171.970 51.060 -171.950 ;
        RECT 148.140 -246.490 150.450 -144.220 ;
        RECT 147.590 -249.330 151.420 -246.490 ;
      LAYER via ;
        RECT -194.640 -121.020 -193.900 -120.530 ;
        RECT 148.800 -248.330 149.970 -247.510 ;
      LAYER met2 ;
        RECT -340.150 -298.900 -330.150 276.100 ;
        RECT -195.720 -298.890 -192.870 -119.590 ;
        RECT 147.840 -249.070 151.070 -246.810 ;
        RECT 148.400 -298.690 150.580 -249.070 ;
        RECT 179.850 -298.900 189.850 276.100 ;
      LAYER via2 ;
        RECT -337.650 268.600 -332.650 273.600 ;
        RECT 182.350 268.600 187.350 273.600 ;
        RECT -337.650 -296.400 -332.650 -291.400 ;
        RECT -194.760 -297.790 -193.910 -289.600 ;
        RECT 148.820 -297.540 149.670 -289.580 ;
        RECT 182.350 -296.400 187.350 -291.400 ;
      LAYER met3 ;
        RECT -400.150 266.100 249.850 276.100 ;
        RECT -400.150 -298.900 249.850 -288.900 ;
    END
  END vdda1
  PIN vssd1
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 41.130 209.990 44.230 212.100 ;
        RECT 42.160 198.600 45.260 200.710 ;
        RECT 42.050 195.140 45.150 197.250 ;
        RECT 42.030 190.230 45.130 192.340 ;
        RECT 42.320 178.310 45.420 180.420 ;
        RECT 42.210 174.850 45.310 176.960 ;
        RECT 42.190 169.940 45.290 172.050 ;
        RECT -6.910 148.570 -3.810 150.680 ;
        RECT 71.020 148.140 74.120 150.250 ;
        RECT -12.670 141.330 9.910 144.110 ;
        RECT 65.260 140.900 87.840 143.680 ;
        RECT -12.670 135.460 9.910 138.240 ;
        RECT 65.260 135.030 87.840 137.810 ;
        RECT -12.720 129.160 9.860 131.940 ;
        RECT 65.210 128.730 87.790 131.510 ;
        RECT -12.930 123.340 9.650 126.120 ;
        RECT 65.000 122.910 87.580 125.690 ;
        RECT -2.600 81.140 19.980 83.920 ;
        RECT 63.960 82.430 86.540 85.210 ;
        RECT 20.040 42.430 32.850 45.090 ;
        RECT 84.730 44.970 97.540 47.630 ;
        RECT -226.850 30.650 -224.740 33.750 ;
        RECT -220.280 16.930 -217.500 39.510 ;
        RECT -214.410 16.930 -211.630 39.510 ;
        RECT -208.110 16.980 -205.330 39.560 ;
        RECT -202.290 17.190 -199.510 39.770 ;
        RECT 65.810 35.330 88.390 38.110 ;
        RECT 0.990 32.340 23.570 35.120 ;
        RECT -160.090 6.860 -157.310 29.440 ;
        RECT -121.260 -6.010 -118.600 6.800 ;
        RECT -111.290 3.270 -108.510 25.850 ;
        RECT 0.000 0.000 8.020 6.760 ;
        RECT -288.270 -17.390 -286.160 -14.290 ;
        RECT -276.880 -18.420 -274.770 -15.320 ;
        RECT -273.420 -18.310 -271.310 -15.210 ;
        RECT -268.510 -18.290 -266.400 -15.190 ;
        RECT -256.590 -18.580 -254.480 -15.480 ;
        RECT -253.130 -18.470 -251.020 -15.370 ;
        RECT -248.220 -18.450 -246.110 -15.350 ;
        RECT -226.420 -47.280 -224.310 -44.180 ;
        RECT -219.850 -61.000 -217.070 -38.420 ;
        RECT -213.980 -61.000 -211.200 -38.420 ;
        RECT -207.680 -60.950 -204.900 -38.370 ;
        RECT -201.860 -60.740 -199.080 -38.160 ;
        RECT -161.380 -59.700 -158.600 -37.120 ;
        RECT -123.800 -70.700 -121.140 -57.890 ;
        RECT -114.280 -61.550 -111.500 -38.970 ;
        RECT 3.410 -61.010 25.990 -58.230 ;
        RECT 68.230 -64.000 90.810 -61.220 ;
        RECT 22.460 -70.980 35.270 -68.320 ;
        RECT 87.150 -73.520 99.960 -70.860 ;
        RECT -0.180 -109.810 22.400 -107.030 ;
        RECT 66.380 -111.100 88.960 -108.320 ;
        RECT -10.510 -152.010 12.070 -149.230 ;
        RECT 67.420 -151.580 90.000 -148.800 ;
        RECT -10.300 -157.830 12.280 -155.050 ;
        RECT 67.630 -157.400 90.210 -154.620 ;
        RECT -10.250 -164.130 12.330 -161.350 ;
        RECT 67.680 -163.700 90.260 -160.920 ;
        RECT -10.250 -170.000 12.330 -167.220 ;
        RECT 67.680 -169.570 90.260 -166.790 ;
        RECT -4.490 -176.570 -1.390 -174.460 ;
        RECT 73.440 -176.140 76.540 -174.030 ;
        RECT 44.610 -197.940 47.710 -195.830 ;
        RECT 44.630 -202.850 47.730 -200.740 ;
        RECT 44.740 -206.310 47.840 -204.200 ;
        RECT 44.450 -218.230 47.550 -216.120 ;
        RECT 44.470 -223.140 47.570 -221.030 ;
        RECT 44.580 -226.600 47.680 -224.490 ;
        RECT 43.550 -237.990 46.650 -235.880 ;
      LAYER li1 ;
        RECT 41.310 211.750 44.050 211.920 ;
        RECT 41.310 210.340 41.480 211.750 ;
        RECT 42.160 211.180 43.200 211.350 ;
        RECT 43.880 210.340 44.050 211.750 ;
        RECT 41.310 210.170 44.050 210.340 ;
        RECT 42.340 200.360 45.080 200.530 ;
        RECT 42.340 198.950 42.510 200.360 ;
        RECT 44.910 198.950 45.080 200.360 ;
        RECT 42.340 198.780 45.080 198.950 ;
        RECT 42.230 196.900 44.970 197.070 ;
        RECT 42.230 195.490 42.400 196.900 ;
        RECT 43.080 195.890 44.120 196.060 ;
        RECT 43.830 195.490 44.030 195.500 ;
        RECT 44.800 195.490 44.970 196.900 ;
        RECT 42.230 195.320 44.970 195.490 ;
        RECT 42.210 191.990 44.950 192.160 ;
        RECT 42.210 190.580 42.380 191.990 ;
        RECT 43.060 191.420 44.100 191.590 ;
        RECT 44.780 190.580 44.950 191.990 ;
        RECT 42.210 190.410 44.950 190.580 ;
        RECT 42.500 180.070 45.240 180.240 ;
        RECT 42.500 178.660 42.670 180.070 ;
        RECT 45.070 178.660 45.240 180.070 ;
        RECT 42.500 178.490 45.240 178.660 ;
        RECT 42.390 176.610 45.130 176.780 ;
        RECT 42.390 175.200 42.560 176.610 ;
        RECT 43.240 175.600 44.280 175.770 ;
        RECT 43.990 175.200 44.190 175.210 ;
        RECT 44.960 175.200 45.130 176.610 ;
        RECT 42.390 175.030 45.130 175.200 ;
        RECT 42.370 171.700 45.110 171.870 ;
        RECT 42.370 170.290 42.540 171.700 ;
        RECT 43.220 171.130 44.260 171.300 ;
        RECT 44.940 170.290 45.110 171.700 ;
        RECT 42.370 170.120 45.110 170.290 ;
        RECT -5.790 150.500 -4.910 150.510 ;
        RECT -6.730 150.330 -3.990 150.500 ;
        RECT -6.730 148.920 -6.560 150.330 ;
        RECT -5.790 149.930 -4.910 150.330 ;
        RECT -5.880 149.760 -4.840 149.930 ;
        RECT -4.160 148.920 -3.990 150.330 ;
        RECT 72.140 150.070 73.020 150.080 ;
        RECT -6.730 148.750 -3.990 148.920 ;
        RECT 71.200 149.900 73.940 150.070 ;
        RECT 71.200 148.490 71.370 149.900 ;
        RECT 72.140 149.500 73.020 149.900 ;
        RECT 72.050 149.330 73.090 149.500 ;
        RECT 73.770 148.490 73.940 149.900 ;
        RECT 71.200 148.320 73.940 148.490 ;
        RECT -12.430 143.700 9.670 143.870 ;
        RECT -12.430 143.390 -12.260 143.700 ;
        RECT -12.430 142.050 -12.250 143.390 ;
        RECT -12.430 141.740 -12.260 142.050 ;
        RECT 9.500 141.740 9.670 143.700 ;
        RECT -12.430 141.570 9.670 141.740 ;
        RECT 65.500 143.270 87.600 143.440 ;
        RECT 65.500 142.960 65.670 143.270 ;
        RECT 65.500 141.620 65.680 142.960 ;
        RECT 65.500 141.310 65.670 141.620 ;
        RECT 87.430 141.310 87.600 143.270 ;
        RECT 65.500 141.140 87.600 141.310 ;
        RECT -12.430 137.830 9.670 138.000 ;
        RECT -12.430 135.870 -12.260 137.830 ;
        RECT -11.400 136.370 8.640 136.540 ;
        RECT 9.500 135.870 9.670 137.830 ;
        RECT -12.430 135.700 9.670 135.870 ;
        RECT 65.500 137.400 87.600 137.570 ;
        RECT 65.500 135.440 65.670 137.400 ;
        RECT 66.530 135.940 86.570 136.110 ;
        RECT 87.430 135.440 87.600 137.400 ;
        RECT 65.500 135.270 87.600 135.440 ;
        RECT -12.480 131.530 9.620 131.700 ;
        RECT -12.480 129.570 -12.310 131.530 ;
        RECT -12.000 131.520 -10.810 131.530 ;
        RECT -11.450 130.860 8.590 131.030 ;
        RECT 9.450 129.570 9.620 131.530 ;
        RECT -12.480 129.400 9.620 129.570 ;
        RECT 65.450 131.100 87.550 131.270 ;
        RECT 65.450 129.140 65.620 131.100 ;
        RECT 65.930 131.090 67.120 131.100 ;
        RECT 66.480 130.430 86.520 130.600 ;
        RECT 87.380 129.140 87.550 131.100 ;
        RECT 65.450 128.970 87.550 129.140 ;
        RECT -12.210 125.880 -10.230 125.900 ;
        RECT -12.690 125.710 9.410 125.880 ;
        RECT -12.690 123.750 -12.520 125.710 ;
        RECT 9.240 123.750 9.410 125.710 ;
        RECT 65.720 125.450 67.700 125.470 ;
        RECT -12.690 123.580 9.410 123.750 ;
        RECT 65.240 125.280 87.340 125.450 ;
        RECT 65.240 123.320 65.410 125.280 ;
        RECT 87.170 123.320 87.340 125.280 ;
        RECT 65.240 123.150 87.340 123.320 ;
        RECT 64.200 84.800 86.300 84.970 ;
        RECT -2.360 83.510 19.740 83.680 ;
        RECT -2.360 81.550 -2.190 83.510 ;
        RECT 19.570 81.550 19.740 83.510 ;
        RECT 64.200 82.840 64.370 84.800 ;
        RECT 86.130 82.840 86.300 84.800 ;
        RECT 64.200 82.670 86.300 82.840 ;
        RECT 65.350 82.660 65.970 82.670 ;
        RECT -2.360 81.380 19.740 81.550 ;
        RECT -1.210 81.370 -0.590 81.380 ;
        RECT 84.910 47.280 97.360 47.450 ;
        RECT 84.910 45.320 85.080 47.280 ;
        RECT 96.460 46.720 96.630 46.800 ;
        RECT 94.645 45.880 96.630 46.720 ;
        RECT 96.460 45.800 96.630 45.880 ;
        RECT 97.190 45.320 97.360 47.280 ;
        RECT 84.910 45.150 97.360 45.320 ;
        RECT 20.220 44.740 32.670 44.910 ;
        RECT 20.220 42.780 20.390 44.740 ;
        RECT 31.770 44.180 31.940 44.260 ;
        RECT 29.955 43.340 31.940 44.180 ;
        RECT 31.770 43.260 31.940 43.340 ;
        RECT 32.500 42.780 32.670 44.740 ;
        RECT 20.220 42.610 32.670 42.780 ;
        RECT -202.050 39.360 -199.750 39.530 ;
        RECT -220.040 39.100 -217.740 39.270 ;
        RECT -226.670 33.400 -224.920 33.570 ;
        RECT -226.670 32.630 -226.500 33.400 ;
        RECT -226.100 32.630 -225.930 32.720 ;
        RECT -226.680 31.750 -225.930 32.630 ;
        RECT -226.670 31.000 -226.500 31.750 ;
        RECT -226.100 31.680 -225.930 31.750 ;
        RECT -225.090 31.000 -224.920 33.400 ;
        RECT -226.670 30.830 -224.920 31.000 ;
        RECT -220.040 17.340 -219.870 39.100 ;
        RECT -219.560 39.090 -218.220 39.100 ;
        RECT -217.910 17.340 -217.740 39.100 ;
        RECT -220.040 17.170 -217.740 17.340 ;
        RECT -214.170 39.100 -211.870 39.270 ;
        RECT -214.170 17.340 -214.000 39.100 ;
        RECT -212.710 18.200 -212.540 38.240 ;
        RECT -212.040 17.340 -211.870 39.100 ;
        RECT -214.170 17.170 -211.870 17.340 ;
        RECT -207.870 39.150 -205.570 39.320 ;
        RECT -207.870 38.840 -207.700 39.150 ;
        RECT -207.870 37.650 -207.690 38.840 ;
        RECT -207.870 17.390 -207.700 37.650 ;
        RECT -207.200 18.250 -207.030 38.290 ;
        RECT -205.740 17.390 -205.570 39.150 ;
        RECT -202.050 39.050 -201.880 39.360 ;
        RECT -202.070 37.070 -201.880 39.050 ;
        RECT -202.050 17.600 -201.880 37.070 ;
        RECT -199.920 17.600 -199.750 39.360 ;
        RECT 66.050 37.700 88.150 37.870 ;
        RECT 66.050 35.740 66.220 37.700 ;
        RECT 87.980 35.740 88.150 37.700 ;
        RECT 66.050 35.570 88.150 35.740 ;
        RECT 67.200 35.560 67.820 35.570 ;
        RECT 1.230 34.710 23.330 34.880 ;
        RECT 1.230 32.750 1.400 34.710 ;
        RECT 23.160 32.750 23.330 34.710 ;
        RECT 1.230 32.580 23.330 32.750 ;
        RECT 2.380 32.570 3.000 32.580 ;
        RECT -202.050 17.430 -199.750 17.600 ;
        RECT -159.850 29.030 -157.550 29.200 ;
        RECT -207.870 17.220 -205.570 17.390 ;
        RECT -159.850 7.270 -159.680 29.030 ;
        RECT -157.720 28.050 -157.550 29.030 ;
        RECT -157.720 27.430 -157.540 28.050 ;
        RECT -157.720 7.270 -157.550 27.430 ;
        RECT -159.850 7.100 -157.550 7.270 ;
        RECT -111.050 25.440 -108.750 25.610 ;
        RECT -121.080 6.450 -118.780 6.620 ;
        RECT -121.080 -5.660 -120.910 6.450 ;
        RECT -120.350 -4.930 -119.510 -3.115 ;
        RECT -120.430 -5.100 -119.430 -4.930 ;
        RECT -118.950 -5.660 -118.780 6.450 ;
        RECT -111.050 3.680 -110.880 25.440 ;
        RECT -108.920 24.460 -108.750 25.440 ;
        RECT -108.920 23.840 -108.740 24.460 ;
        RECT -108.920 3.680 -108.750 23.840 ;
        RECT 0.440 4.640 1.040 5.640 ;
        RECT 4.520 4.660 5.120 5.660 ;
        RECT -111.050 3.510 -108.750 3.680 ;
        RECT 0.400 1.200 1.000 2.200 ;
        RECT 4.460 1.220 5.060 2.220 ;
        RECT -121.080 -5.830 -118.780 -5.660 ;
        RECT -288.090 -14.640 -286.340 -14.470 ;
        RECT -288.090 -17.040 -287.920 -14.640 ;
        RECT -287.520 -16.360 -287.350 -15.320 ;
        RECT -286.510 -17.040 -286.340 -14.640 ;
        RECT -288.090 -17.210 -286.340 -17.040 ;
        RECT -276.700 -15.670 -274.950 -15.500 ;
        RECT -276.700 -18.070 -276.530 -15.670 ;
        RECT -275.120 -18.070 -274.950 -15.670 ;
        RECT -276.700 -18.240 -274.950 -18.070 ;
        RECT -273.240 -15.560 -271.490 -15.390 ;
        RECT -273.240 -17.960 -273.070 -15.560 ;
        RECT -272.230 -17.280 -272.060 -16.240 ;
        RECT -271.660 -16.990 -271.490 -15.560 ;
        RECT -271.670 -17.190 -271.490 -16.990 ;
        RECT -271.660 -17.960 -271.490 -17.190 ;
        RECT -273.240 -18.130 -271.490 -17.960 ;
        RECT -268.330 -15.540 -266.580 -15.370 ;
        RECT -268.330 -17.940 -268.160 -15.540 ;
        RECT -267.760 -17.260 -267.590 -16.220 ;
        RECT -266.750 -17.940 -266.580 -15.540 ;
        RECT -268.330 -18.110 -266.580 -17.940 ;
        RECT -256.410 -15.830 -254.660 -15.660 ;
        RECT -256.410 -18.230 -256.240 -15.830 ;
        RECT -254.830 -18.230 -254.660 -15.830 ;
        RECT -256.410 -18.400 -254.660 -18.230 ;
        RECT -252.950 -15.720 -251.200 -15.550 ;
        RECT -252.950 -18.120 -252.780 -15.720 ;
        RECT -251.940 -17.440 -251.770 -16.400 ;
        RECT -251.370 -17.150 -251.200 -15.720 ;
        RECT -251.380 -17.350 -251.200 -17.150 ;
        RECT -251.370 -18.120 -251.200 -17.350 ;
        RECT -252.950 -18.290 -251.200 -18.120 ;
        RECT -248.040 -15.700 -246.290 -15.530 ;
        RECT -248.040 -18.100 -247.870 -15.700 ;
        RECT -247.470 -17.420 -247.300 -16.380 ;
        RECT -246.460 -18.100 -246.290 -15.700 ;
        RECT -248.040 -18.270 -246.290 -18.100 ;
        RECT -161.140 -37.530 -158.840 -37.360 ;
        RECT -201.620 -38.570 -199.320 -38.400 ;
        RECT -219.610 -38.830 -217.310 -38.660 ;
        RECT -226.240 -44.530 -224.490 -44.360 ;
        RECT -226.240 -45.300 -226.070 -44.530 ;
        RECT -225.670 -45.300 -225.500 -45.210 ;
        RECT -226.250 -46.180 -225.500 -45.300 ;
        RECT -226.240 -46.930 -226.070 -46.180 ;
        RECT -225.670 -46.250 -225.500 -46.180 ;
        RECT -224.660 -46.930 -224.490 -44.530 ;
        RECT -226.240 -47.100 -224.490 -46.930 ;
        RECT -219.610 -60.590 -219.440 -38.830 ;
        RECT -219.130 -38.840 -217.790 -38.830 ;
        RECT -217.480 -60.590 -217.310 -38.830 ;
        RECT -219.610 -60.760 -217.310 -60.590 ;
        RECT -213.740 -38.830 -211.440 -38.660 ;
        RECT -213.740 -60.590 -213.570 -38.830 ;
        RECT -212.280 -59.730 -212.110 -39.690 ;
        RECT -211.610 -60.590 -211.440 -38.830 ;
        RECT -213.740 -60.760 -211.440 -60.590 ;
        RECT -207.440 -38.780 -205.140 -38.610 ;
        RECT -207.440 -39.090 -207.270 -38.780 ;
        RECT -207.440 -40.280 -207.260 -39.090 ;
        RECT -207.440 -60.540 -207.270 -40.280 ;
        RECT -206.770 -59.680 -206.600 -39.640 ;
        RECT -205.310 -60.540 -205.140 -38.780 ;
        RECT -201.620 -38.880 -201.450 -38.570 ;
        RECT -201.640 -40.860 -201.450 -38.880 ;
        RECT -201.620 -60.330 -201.450 -40.860 ;
        RECT -199.490 -60.330 -199.320 -38.570 ;
        RECT -161.140 -59.290 -160.970 -37.530 ;
        RECT -159.010 -38.510 -158.840 -37.530 ;
        RECT -159.010 -39.130 -158.830 -38.510 ;
        RECT -159.010 -59.290 -158.840 -39.130 ;
        RECT -114.040 -39.380 -111.740 -39.210 ;
        RECT -161.140 -59.460 -158.840 -59.290 ;
        RECT -123.620 -58.240 -121.320 -58.070 ;
        RECT -201.620 -60.500 -199.320 -60.330 ;
        RECT -207.440 -60.710 -205.140 -60.540 ;
        RECT -123.620 -70.350 -123.450 -58.240 ;
        RECT -122.890 -69.620 -122.050 -67.805 ;
        RECT -122.970 -69.790 -121.970 -69.620 ;
        RECT -121.490 -70.350 -121.320 -58.240 ;
        RECT -114.040 -61.140 -113.870 -39.380 ;
        RECT -111.910 -40.360 -111.740 -39.380 ;
        RECT -111.910 -40.980 -111.730 -40.360 ;
        RECT -111.910 -61.140 -111.740 -40.980 ;
        RECT 4.800 -58.470 5.420 -58.460 ;
        RECT 3.650 -58.640 25.750 -58.470 ;
        RECT 3.650 -60.600 3.820 -58.640 ;
        RECT 25.580 -60.600 25.750 -58.640 ;
        RECT 3.650 -60.770 25.750 -60.600 ;
        RECT -114.040 -61.310 -111.740 -61.140 ;
        RECT 69.620 -61.460 70.240 -61.450 ;
        RECT 68.470 -61.630 90.570 -61.460 ;
        RECT 68.470 -63.590 68.640 -61.630 ;
        RECT 90.400 -63.590 90.570 -61.630 ;
        RECT 68.470 -63.760 90.570 -63.590 ;
        RECT -123.620 -70.520 -121.320 -70.350 ;
        RECT 22.640 -68.670 35.090 -68.500 ;
        RECT 22.640 -70.630 22.810 -68.670 ;
        RECT 34.190 -69.230 34.360 -69.150 ;
        RECT 32.375 -70.070 34.360 -69.230 ;
        RECT 34.190 -70.150 34.360 -70.070 ;
        RECT 34.920 -70.630 35.090 -68.670 ;
        RECT 22.640 -70.800 35.090 -70.630 ;
        RECT 87.330 -71.210 99.780 -71.040 ;
        RECT 87.330 -73.170 87.500 -71.210 ;
        RECT 98.880 -71.770 99.050 -71.690 ;
        RECT 97.065 -72.610 99.050 -71.770 ;
        RECT 98.880 -72.690 99.050 -72.610 ;
        RECT 99.610 -73.170 99.780 -71.210 ;
        RECT 87.330 -73.340 99.780 -73.170 ;
        RECT 1.210 -107.270 1.830 -107.260 ;
        RECT 0.060 -107.440 22.160 -107.270 ;
        RECT 0.060 -109.400 0.230 -107.440 ;
        RECT 21.990 -109.400 22.160 -107.440 ;
        RECT 67.770 -108.560 68.390 -108.550 ;
        RECT 0.060 -109.570 22.160 -109.400 ;
        RECT 66.620 -108.730 88.720 -108.560 ;
        RECT 66.620 -110.690 66.790 -108.730 ;
        RECT 88.550 -110.690 88.720 -108.730 ;
        RECT 66.620 -110.860 88.720 -110.690 ;
        RECT 67.660 -149.210 89.760 -149.040 ;
        RECT -10.270 -149.640 11.830 -149.470 ;
        RECT -10.270 -151.600 -10.100 -149.640 ;
        RECT 11.660 -151.600 11.830 -149.640 ;
        RECT 67.660 -151.170 67.830 -149.210 ;
        RECT 89.590 -151.170 89.760 -149.210 ;
        RECT 67.660 -151.340 89.760 -151.170 ;
        RECT 68.140 -151.360 70.120 -151.340 ;
        RECT -10.270 -151.770 11.830 -151.600 ;
        RECT -9.790 -151.790 -7.810 -151.770 ;
        RECT 67.870 -155.030 89.970 -154.860 ;
        RECT -10.060 -155.460 12.040 -155.290 ;
        RECT -10.060 -157.420 -9.890 -155.460 ;
        RECT -9.030 -156.920 11.010 -156.750 ;
        RECT -9.580 -157.420 -8.390 -157.410 ;
        RECT 11.870 -157.420 12.040 -155.460 ;
        RECT 67.870 -156.990 68.040 -155.030 ;
        RECT 68.900 -156.490 88.940 -156.320 ;
        RECT 68.350 -156.990 69.540 -156.980 ;
        RECT 89.800 -156.990 89.970 -155.030 ;
        RECT 67.870 -157.160 89.970 -156.990 ;
        RECT -10.060 -157.590 12.040 -157.420 ;
        RECT 67.920 -161.330 90.020 -161.160 ;
        RECT -10.010 -161.760 12.090 -161.590 ;
        RECT -10.010 -163.720 -9.840 -161.760 ;
        RECT -8.980 -162.430 11.060 -162.260 ;
        RECT 11.920 -163.720 12.090 -161.760 ;
        RECT 67.920 -163.290 68.090 -161.330 ;
        RECT 68.950 -162.000 88.990 -161.830 ;
        RECT 89.850 -163.290 90.020 -161.330 ;
        RECT 67.920 -163.460 90.020 -163.290 ;
        RECT -10.010 -163.890 12.090 -163.720 ;
        RECT 67.920 -167.200 90.020 -167.030 ;
        RECT -10.010 -167.630 12.090 -167.460 ;
        RECT -10.010 -167.940 -9.840 -167.630 ;
        RECT -10.010 -169.280 -9.830 -167.940 ;
        RECT -10.010 -169.590 -9.840 -169.280 ;
        RECT 11.920 -169.590 12.090 -167.630 ;
        RECT 67.920 -167.510 68.090 -167.200 ;
        RECT 67.920 -168.850 68.100 -167.510 ;
        RECT 67.920 -169.160 68.090 -168.850 ;
        RECT 89.850 -169.160 90.020 -167.200 ;
        RECT 67.920 -169.330 90.020 -169.160 ;
        RECT -10.010 -169.760 12.090 -169.590 ;
        RECT 73.620 -174.380 76.360 -174.210 ;
        RECT -4.310 -174.810 -1.570 -174.640 ;
        RECT -4.310 -176.220 -4.140 -174.810 ;
        RECT -3.460 -175.820 -2.420 -175.650 ;
        RECT -3.370 -176.220 -2.490 -175.820 ;
        RECT -1.740 -176.220 -1.570 -174.810 ;
        RECT 73.620 -175.790 73.790 -174.380 ;
        RECT 74.470 -175.390 75.510 -175.220 ;
        RECT 74.560 -175.790 75.440 -175.390 ;
        RECT 76.190 -175.790 76.360 -174.380 ;
        RECT 73.620 -175.960 76.360 -175.790 ;
        RECT 74.560 -175.970 75.440 -175.960 ;
        RECT -4.310 -176.390 -1.570 -176.220 ;
        RECT -3.370 -176.400 -2.490 -176.390 ;
        RECT 44.790 -196.180 47.530 -196.010 ;
        RECT 44.790 -197.590 44.960 -196.180 ;
        RECT 45.640 -197.190 46.680 -197.020 ;
        RECT 47.360 -197.590 47.530 -196.180 ;
        RECT 44.790 -197.760 47.530 -197.590 ;
        RECT 44.810 -201.090 47.550 -200.920 ;
        RECT 44.810 -202.500 44.980 -201.090 ;
        RECT 46.410 -201.100 46.610 -201.090 ;
        RECT 45.660 -201.660 46.700 -201.490 ;
        RECT 47.380 -202.500 47.550 -201.090 ;
        RECT 44.810 -202.670 47.550 -202.500 ;
        RECT 44.920 -204.550 47.660 -204.380 ;
        RECT 44.920 -205.960 45.090 -204.550 ;
        RECT 47.490 -205.960 47.660 -204.550 ;
        RECT 44.920 -206.130 47.660 -205.960 ;
        RECT 44.630 -216.470 47.370 -216.300 ;
        RECT 44.630 -217.880 44.800 -216.470 ;
        RECT 45.480 -217.480 46.520 -217.310 ;
        RECT 47.200 -217.880 47.370 -216.470 ;
        RECT 44.630 -218.050 47.370 -217.880 ;
        RECT 44.650 -221.380 47.390 -221.210 ;
        RECT 44.650 -222.790 44.820 -221.380 ;
        RECT 46.250 -221.390 46.450 -221.380 ;
        RECT 45.500 -221.950 46.540 -221.780 ;
        RECT 47.220 -222.790 47.390 -221.380 ;
        RECT 44.650 -222.960 47.390 -222.790 ;
        RECT 44.760 -224.840 47.500 -224.670 ;
        RECT 44.760 -226.250 44.930 -224.840 ;
        RECT 47.330 -226.250 47.500 -224.840 ;
        RECT 44.760 -226.420 47.500 -226.250 ;
        RECT 43.730 -236.230 46.470 -236.060 ;
        RECT 43.730 -237.640 43.900 -236.230 ;
        RECT 44.580 -237.240 45.620 -237.070 ;
        RECT 46.300 -237.640 46.470 -236.230 ;
        RECT 43.730 -237.810 46.470 -237.640 ;
      LAYER mcon ;
        RECT 42.850 211.750 43.120 211.920 ;
        RECT 42.240 211.180 43.120 211.350 ;
        RECT 42.340 199.260 42.510 200.050 ;
        RECT 42.230 195.800 42.400 196.590 ;
        RECT 43.160 195.890 44.040 196.060 ;
        RECT 43.830 195.320 44.030 195.500 ;
        RECT 43.760 191.990 44.010 192.160 ;
        RECT 43.140 191.420 44.020 191.590 ;
        RECT 42.500 178.970 42.670 179.760 ;
        RECT 42.390 175.510 42.560 176.300 ;
        RECT 43.320 175.600 44.200 175.770 ;
        RECT 43.990 175.030 44.190 175.210 ;
        RECT 43.920 171.700 44.170 171.870 ;
        RECT 43.300 171.130 44.180 171.300 ;
        RECT -5.800 149.760 -4.920 149.930 ;
        RECT -6.250 148.750 -4.470 148.920 ;
        RECT 72.130 149.330 73.010 149.500 ;
        RECT 71.680 148.320 73.460 148.490 ;
        RECT -12.430 142.050 -12.250 143.390 ;
        RECT 65.500 141.620 65.680 142.960 ;
        RECT -11.320 136.370 8.560 136.540 ;
        RECT -11.950 135.700 -10.760 135.870 ;
        RECT -3.680 135.700 -2.740 135.870 ;
        RECT 7.690 135.700 9.190 135.870 ;
        RECT 66.610 135.940 86.490 136.110 ;
        RECT 65.980 135.270 67.170 135.440 ;
        RECT 74.250 135.270 75.190 135.440 ;
        RECT 85.620 135.270 87.120 135.440 ;
        RECT -11.370 130.860 8.510 131.030 ;
        RECT 66.560 130.430 86.440 130.600 ;
        RECT -12.210 125.710 -10.230 125.900 ;
        RECT 65.720 125.280 67.700 125.470 ;
        RECT 94.645 45.880 96.630 46.720 ;
        RECT 29.955 43.340 31.940 44.180 ;
        RECT -226.100 31.760 -225.930 32.640 ;
        RECT -225.090 31.310 -224.920 33.090 ;
        RECT -212.710 18.280 -212.540 38.160 ;
        RECT -212.040 37.600 -211.870 38.790 ;
        RECT -212.040 29.580 -211.870 30.520 ;
        RECT -212.040 17.650 -211.870 19.150 ;
        RECT -207.860 37.650 -207.690 38.840 ;
        RECT -207.200 18.330 -207.030 38.210 ;
        RECT -202.070 37.070 -201.880 39.050 ;
        RECT -157.720 27.430 -157.540 28.050 ;
        RECT -120.350 -5.100 -119.510 -3.115 ;
        RECT -108.920 23.840 -108.740 24.460 ;
        RECT 0.540 4.735 0.940 5.540 ;
        RECT 4.620 4.755 5.020 5.560 ;
        RECT 0.500 1.295 0.900 2.100 ;
        RECT 4.560 1.315 4.960 2.120 ;
        RECT -288.090 -16.280 -287.920 -16.010 ;
        RECT -287.520 -16.280 -287.350 -15.400 ;
        RECT -276.220 -15.670 -275.430 -15.500 ;
        RECT -272.760 -15.560 -271.970 -15.390 ;
        RECT -272.230 -17.200 -272.060 -16.320 ;
        RECT -271.670 -17.190 -271.490 -16.990 ;
        RECT -268.330 -17.170 -268.160 -16.920 ;
        RECT -267.760 -17.180 -267.590 -16.300 ;
        RECT -255.930 -15.830 -255.140 -15.660 ;
        RECT -252.470 -15.720 -251.680 -15.550 ;
        RECT -251.940 -17.360 -251.770 -16.480 ;
        RECT -251.380 -17.350 -251.200 -17.150 ;
        RECT -248.040 -17.330 -247.870 -17.080 ;
        RECT -247.470 -17.340 -247.300 -16.460 ;
        RECT -225.670 -46.170 -225.500 -45.290 ;
        RECT -224.660 -46.620 -224.490 -44.840 ;
        RECT -212.280 -59.650 -212.110 -39.770 ;
        RECT -211.610 -40.330 -211.440 -39.140 ;
        RECT -211.610 -48.350 -211.440 -47.410 ;
        RECT -211.610 -60.280 -211.440 -58.780 ;
        RECT -207.430 -40.280 -207.260 -39.090 ;
        RECT -206.770 -59.600 -206.600 -39.720 ;
        RECT -201.640 -40.860 -201.450 -38.880 ;
        RECT -159.010 -39.130 -158.830 -38.510 ;
        RECT -122.890 -69.790 -122.050 -67.805 ;
        RECT -111.910 -40.980 -111.730 -40.360 ;
        RECT 4.800 -58.640 5.420 -58.460 ;
        RECT 69.620 -61.630 70.240 -61.450 ;
        RECT 32.375 -70.070 34.360 -69.230 ;
        RECT 97.065 -72.610 99.050 -71.770 ;
        RECT 1.210 -107.440 1.830 -107.260 ;
        RECT 67.770 -108.730 68.390 -108.550 ;
        RECT -8.950 -156.920 10.930 -156.750 ;
        RECT -9.580 -157.580 -8.390 -157.410 ;
        RECT 68.980 -156.490 88.860 -156.320 ;
        RECT 68.350 -157.150 69.540 -156.980 ;
        RECT 68.400 -161.330 69.590 -161.160 ;
        RECT 76.670 -161.330 77.610 -161.160 ;
        RECT 88.040 -161.330 89.540 -161.160 ;
        RECT -9.530 -161.760 -8.340 -161.590 ;
        RECT -1.260 -161.760 -0.320 -161.590 ;
        RECT 10.110 -161.760 11.610 -161.590 ;
        RECT -8.900 -162.430 10.980 -162.260 ;
        RECT 69.030 -162.000 88.910 -161.830 ;
        RECT -10.010 -169.280 -9.830 -167.940 ;
        RECT 67.920 -168.850 68.100 -167.510 ;
        RECT 74.100 -174.380 75.880 -174.210 ;
        RECT -3.830 -174.810 -2.050 -174.640 ;
        RECT -3.380 -175.820 -2.500 -175.650 ;
        RECT 74.550 -175.390 75.430 -175.220 ;
        RECT 45.720 -197.190 46.600 -197.020 ;
        RECT 46.340 -197.760 46.590 -197.590 ;
        RECT 44.810 -202.190 44.980 -201.400 ;
        RECT 45.740 -201.660 46.620 -201.490 ;
        RECT 44.920 -205.650 45.090 -204.860 ;
        RECT 45.560 -217.480 46.440 -217.310 ;
        RECT 46.180 -218.050 46.430 -217.880 ;
        RECT 44.650 -222.480 44.820 -221.690 ;
        RECT 45.580 -221.950 46.460 -221.780 ;
        RECT 44.760 -225.940 44.930 -225.150 ;
        RECT 44.660 -237.240 45.540 -237.070 ;
        RECT 45.270 -237.810 45.540 -237.640 ;
      LAYER met1 ;
        RECT 39.990 211.680 43.190 212.010 ;
        RECT 39.990 211.630 43.150 211.680 ;
        RECT 39.990 198.320 40.270 211.630 ;
        RECT 42.850 211.380 43.100 211.630 ;
        RECT 42.180 211.150 43.180 211.380 ;
        RECT 42.280 200.100 42.590 200.140 ;
        RECT 39.680 198.210 40.270 198.320 ;
        RECT 40.930 200.010 41.250 200.050 ;
        RECT 42.270 200.010 42.590 200.100 ;
        RECT 40.930 199.430 42.590 200.010 ;
        RECT 40.930 198.210 41.250 199.430 ;
        RECT 42.270 199.240 42.590 199.430 ;
        RECT 42.280 199.200 42.590 199.240 ;
        RECT 39.590 197.700 41.250 198.210 ;
        RECT -100.030 69.730 -95.810 73.160 ;
        RECT -39.670 72.520 -37.420 146.720 ;
        RECT -32.920 146.630 -31.480 179.470 ;
        RECT -31.220 179.130 9.580 179.230 ;
        RECT -31.220 179.050 37.330 179.130 ;
        RECT 39.680 179.050 40.230 197.700 ;
        RECT 40.930 196.410 41.250 197.700 ;
        RECT 42.100 196.410 42.470 196.680 ;
        RECT 40.930 195.900 42.470 196.410 ;
        RECT 43.110 196.090 44.090 196.110 ;
        RECT 40.930 195.870 41.550 195.900 ;
        RECT 41.090 193.140 41.550 195.870 ;
        RECT 42.100 195.690 42.470 195.900 ;
        RECT 43.100 195.860 44.100 196.090 ;
        RECT 43.110 195.830 44.090 195.860 ;
        RECT 43.840 195.610 44.040 195.830 ;
        RECT 43.720 195.200 44.100 195.610 ;
        RECT 41.090 192.740 44.110 193.140 ;
        RECT 41.090 192.710 41.550 192.740 ;
        RECT 43.800 192.240 44.070 192.740 ;
        RECT 43.680 191.910 44.090 192.240 ;
        RECT 43.740 191.620 44.010 191.910 ;
        RECT 43.080 191.390 44.080 191.620 ;
        RECT 42.440 179.810 42.750 179.850 ;
        RECT -31.220 178.380 40.230 179.050 ;
        RECT -3.470 178.280 40.230 178.380 ;
        RECT 37.070 178.110 40.230 178.280 ;
        RECT 39.680 177.920 40.230 178.110 ;
        RECT 41.090 179.720 41.410 179.760 ;
        RECT 42.430 179.720 42.750 179.810 ;
        RECT 41.090 179.140 42.750 179.720 ;
        RECT 41.090 177.920 41.410 179.140 ;
        RECT 42.430 178.950 42.750 179.140 ;
        RECT 42.440 178.910 42.750 178.950 ;
        RECT 39.680 177.410 41.410 177.920 ;
        RECT 41.090 176.120 41.410 177.410 ;
        RECT 42.260 176.120 42.630 176.390 ;
        RECT 41.090 175.610 42.630 176.120 ;
        RECT 43.270 175.800 44.250 175.820 ;
        RECT 41.090 175.580 41.710 175.610 ;
        RECT 41.250 172.850 41.710 175.580 ;
        RECT 42.260 175.400 42.630 175.610 ;
        RECT 43.260 175.570 44.260 175.800 ;
        RECT 43.270 175.540 44.250 175.570 ;
        RECT 44.000 175.320 44.200 175.540 ;
        RECT 43.880 174.910 44.260 175.320 ;
        RECT 41.250 172.450 44.270 172.850 ;
        RECT 41.250 172.420 41.710 172.450 ;
        RECT 43.960 171.950 44.230 172.450 ;
        RECT 43.840 171.620 44.250 171.950 ;
        RECT 43.900 171.330 44.170 171.620 ;
        RECT 43.240 171.100 44.240 171.330 ;
        RECT -5.870 149.710 -4.860 150.070 ;
        RECT 72.060 149.280 73.070 149.640 ;
        RECT -6.310 148.980 -6.160 149.040 ;
        RECT -37.170 144.620 -31.480 146.630 ;
        RECT -32.920 125.610 -31.480 144.620 ;
        RECT -13.450 148.680 -3.770 148.980 ;
        RECT -13.450 148.640 -6.150 148.680 ;
        RECT -13.450 142.420 -13.290 148.640 ;
        RECT 71.620 148.550 71.770 148.610 ;
        RECT 64.480 148.250 74.160 148.550 ;
        RECT 64.480 148.210 71.780 148.250 ;
        RECT -12.490 142.420 -12.190 143.420 ;
        RECT -13.490 142.050 -12.190 142.420 ;
        RECT -13.460 135.900 -13.240 142.050 ;
        RECT -12.490 141.980 -12.190 142.050 ;
        RECT 64.480 141.990 64.640 148.210 ;
        RECT 65.440 141.990 65.740 142.990 ;
        RECT 64.440 141.620 65.740 141.990 ;
        RECT -11.380 136.340 8.620 136.570 ;
        RECT -11.320 135.930 -10.760 136.340 ;
        RECT -3.680 135.940 -2.740 136.340 ;
        RECT -3.760 135.930 -2.740 135.940 ;
        RECT 7.690 135.930 8.510 136.340 ;
        RECT -13.490 135.890 -13.190 135.900 ;
        RECT -12.000 135.890 -10.670 135.930 ;
        RECT -13.490 135.660 -10.660 135.890 ;
        RECT -13.490 129.440 -13.190 135.660 ;
        RECT -12.000 135.640 -10.670 135.660 ;
        RECT -3.760 135.640 -2.640 135.930 ;
        RECT 7.590 135.640 9.240 135.930 ;
        RECT -11.320 135.630 -10.670 135.640 ;
        RECT -11.320 131.790 -10.760 135.630 ;
        RECT -12.030 131.460 -10.760 131.790 ;
        RECT -11.320 131.060 -10.760 131.460 ;
        RECT -3.680 131.060 -2.740 135.640 ;
        RECT 7.590 135.630 8.510 135.640 ;
        RECT 7.690 131.060 8.510 135.630 ;
        RECT 64.470 135.470 64.690 141.620 ;
        RECT 65.440 141.550 65.740 141.620 ;
        RECT 66.550 135.910 86.550 136.140 ;
        RECT 66.610 135.500 67.170 135.910 ;
        RECT 74.250 135.510 75.190 135.910 ;
        RECT 74.170 135.500 75.190 135.510 ;
        RECT 85.620 135.500 86.440 135.910 ;
        RECT 64.440 135.460 64.740 135.470 ;
        RECT 65.930 135.460 67.260 135.500 ;
        RECT 64.440 135.230 67.270 135.460 ;
        RECT -11.430 130.830 8.570 131.060 ;
        RECT -14.810 127.550 -13.190 129.440 ;
        RECT 64.440 128.360 64.740 135.230 ;
        RECT 65.930 135.210 67.260 135.230 ;
        RECT 74.170 135.210 75.290 135.500 ;
        RECT 85.520 135.210 87.170 135.500 ;
        RECT 66.610 135.200 67.260 135.210 ;
        RECT 66.610 131.360 67.170 135.200 ;
        RECT 65.900 131.030 67.170 131.360 ;
        RECT 66.610 130.630 67.170 131.030 ;
        RECT 74.250 130.630 75.190 135.210 ;
        RECT 85.520 135.200 86.440 135.210 ;
        RECT 85.620 130.630 86.440 135.200 ;
        RECT 66.500 130.400 86.500 130.630 ;
        RECT -13.490 125.980 -13.190 127.550 ;
        RECT 63.750 126.850 64.740 128.360 ;
        RECT -13.490 125.680 -10.170 125.980 ;
        RECT -33.850 124.220 -31.470 125.610 ;
        RECT 64.440 125.550 64.740 126.850 ;
        RECT 64.440 125.250 67.760 125.550 ;
        RECT -33.750 114.670 -32.910 124.220 ;
        RECT -34.690 109.830 -31.880 114.670 ;
        RECT 65.300 82.600 66.020 82.910 ;
        RECT 65.380 82.010 65.970 82.600 ;
        RECT -1.260 81.310 -0.540 81.620 ;
        RECT -1.180 81.010 -0.590 81.310 ;
        RECT -1.270 80.720 -0.590 81.010 ;
        RECT -15.140 72.620 -10.170 73.830 ;
        RECT -26.100 72.520 -10.170 72.620 ;
        RECT -39.670 70.140 -10.170 72.520 ;
        RECT -39.670 70.040 -24.300 70.140 ;
        RECT -99.110 66.750 -97.540 69.730 ;
        RECT -99.400 66.510 -97.540 66.750 ;
        RECT -222.890 64.260 -96.890 66.510 ;
        RECT -222.800 59.760 -220.790 64.010 ;
        RECT -201.780 60.590 -200.390 60.690 ;
        RECT -190.840 60.590 -186.000 61.530 ;
        RECT -201.780 59.760 -186.000 60.590 ;
        RECT -255.640 59.750 -186.000 59.760 ;
        RECT -255.640 58.320 -200.390 59.750 ;
        RECT -190.840 58.720 -186.000 59.750 ;
        RECT -201.780 58.310 -200.390 58.320 ;
        RECT -255.400 30.310 -254.550 58.060 ;
        RECT -148.690 52.940 -146.210 64.260 ;
        RECT -148.790 51.140 -146.210 52.940 ;
        RECT -148.790 41.980 -146.310 51.140 ;
        RECT -205.610 40.330 -203.720 41.650 ;
        RECT -218.590 40.300 -218.220 40.330 ;
        RECT -212.070 40.300 -201.850 40.330 ;
        RECT -218.590 40.290 -201.850 40.300 ;
        RECT -225.150 40.130 -201.850 40.290 ;
        RECT -225.150 33.150 -224.810 40.130 ;
        RECT -218.590 40.080 -201.850 40.130 ;
        RECT -218.590 39.330 -218.220 40.080 ;
        RECT -212.070 40.030 -201.850 40.080 ;
        RECT -219.590 39.030 -218.150 39.330 ;
        RECT -212.060 38.840 -211.830 40.030 ;
        RECT -225.210 33.000 -224.810 33.150 ;
        RECT -225.150 32.990 -224.810 33.000 ;
        RECT -212.740 38.160 -212.510 38.220 ;
        RECT -212.100 38.160 -211.810 38.840 ;
        RECT -207.960 38.160 -207.630 38.870 ;
        RECT -207.230 38.160 -207.000 38.270 ;
        RECT -212.740 37.600 -207.000 38.160 ;
        RECT -226.240 31.700 -225.880 32.710 ;
        RECT -225.150 30.610 -224.850 32.990 ;
        RECT -212.740 30.520 -212.510 37.600 ;
        RECT -212.100 37.510 -211.800 37.600 ;
        RECT -212.060 37.500 -211.830 37.510 ;
        RECT -212.110 30.520 -211.810 30.600 ;
        RECT -207.230 30.520 -207.000 37.600 ;
        RECT -202.150 37.010 -201.850 40.030 ;
        RECT -150.000 37.010 -144.340 41.980 ;
        RECT -99.400 40.210 -97.850 64.260 ;
        RECT -39.670 40.210 -37.420 70.040 ;
        RECT -15.140 68.170 -10.170 70.140 ;
        RECT -1.270 73.600 -0.830 80.720 ;
        RECT -1.270 67.880 2.250 73.600 ;
        RECT -1.270 65.160 -0.830 67.880 ;
        RECT 65.440 65.460 65.880 82.010 ;
        RECT 65.240 65.160 66.030 65.460 ;
        RECT -1.270 64.730 66.030 65.160 ;
        RECT -1.270 63.750 -0.830 64.730 ;
        RECT 65.240 64.670 66.030 64.730 ;
        RECT 94.585 45.850 96.690 46.750 ;
        RECT 29.895 43.310 32.000 44.210 ;
        RECT -99.400 39.150 -37.420 40.210 ;
        RECT -255.400 17.260 -254.450 30.310 ;
        RECT -212.740 29.580 -207.000 30.520 ;
        RECT -212.740 19.150 -212.510 29.580 ;
        RECT -212.100 29.480 -211.810 29.580 ;
        RECT -212.100 19.150 -211.800 19.250 ;
        RECT -207.230 19.150 -207.000 29.580 ;
        RECT -157.790 28.020 -157.480 28.100 ;
        RECT -157.180 28.020 -139.920 28.110 ;
        RECT -157.790 27.670 -139.920 28.020 ;
        RECT -157.790 27.430 -156.890 27.670 ;
        RECT -157.790 27.380 -157.480 27.430 ;
        RECT -149.770 24.590 -144.050 27.670 ;
        RECT -212.740 18.330 -207.000 19.150 ;
        RECT -212.740 18.220 -212.510 18.330 ;
        RECT -212.100 17.600 -211.810 18.330 ;
        RECT -207.230 18.270 -207.000 18.330 ;
        RECT -255.300 -10.230 -254.450 17.260 ;
        RECT -255.300 -10.490 -254.280 -10.230 ;
        RECT -274.380 -12.840 -273.870 -12.750 ;
        RECT -255.220 -12.840 -254.280 -10.490 ;
        RECT -274.490 -13.150 -253.580 -12.840 ;
        RECT -288.180 -13.390 -253.580 -13.150 ;
        RECT -288.180 -13.430 -273.870 -13.390 ;
        RECT -288.180 -16.010 -287.800 -13.430 ;
        RECT -274.380 -14.090 -273.870 -13.430 ;
        RECT -276.220 -14.250 -272.040 -14.090 ;
        RECT -254.090 -14.250 -253.580 -13.390 ;
        RECT -276.220 -14.410 -268.880 -14.250 ;
        RECT -287.550 -16.010 -287.320 -15.340 ;
        RECT -276.180 -15.430 -275.600 -14.410 ;
        RECT -272.580 -14.710 -268.880 -14.410 ;
        RECT -255.930 -14.410 -251.750 -14.250 ;
        RECT -255.930 -14.570 -248.590 -14.410 ;
        RECT -272.580 -15.260 -272.070 -14.710 ;
        RECT -276.270 -15.440 -275.410 -15.430 ;
        RECT -276.310 -15.750 -275.370 -15.440 ;
        RECT -272.850 -15.630 -271.860 -15.260 ;
        RECT -288.180 -16.260 -287.320 -16.010 ;
        RECT -288.180 -16.310 -287.800 -16.260 ;
        RECT -288.180 -16.350 -287.850 -16.310 ;
        RECT -287.550 -16.340 -287.320 -16.260 ;
        RECT -272.260 -16.270 -272.030 -16.260 ;
        RECT -272.280 -17.000 -272.000 -16.270 ;
        RECT -271.780 -17.000 -271.370 -16.880 ;
        RECT -272.280 -17.200 -271.370 -17.000 ;
        RECT -272.280 -17.250 -272.000 -17.200 ;
        RECT -272.260 -17.260 -272.030 -17.250 ;
        RECT -271.780 -17.260 -271.370 -17.200 ;
        RECT -269.310 -16.960 -268.910 -14.710 ;
        RECT -255.890 -15.590 -255.310 -14.570 ;
        RECT -252.290 -14.870 -248.590 -14.570 ;
        RECT -252.290 -15.420 -251.780 -14.870 ;
        RECT -255.980 -15.600 -255.120 -15.590 ;
        RECT -256.020 -15.910 -255.080 -15.600 ;
        RECT -252.560 -15.790 -251.570 -15.420 ;
        RECT -268.410 -16.900 -268.080 -16.840 ;
        RECT -267.790 -16.900 -267.560 -16.240 ;
        RECT -251.970 -16.430 -251.740 -16.420 ;
        RECT -268.410 -16.960 -267.560 -16.900 ;
        RECT -269.310 -17.170 -267.560 -16.960 ;
        RECT -269.310 -17.230 -268.080 -17.170 ;
        RECT -269.310 -17.270 -268.910 -17.230 ;
        RECT -268.410 -17.250 -268.080 -17.230 ;
        RECT -267.790 -17.240 -267.560 -17.170 ;
        RECT -251.990 -17.160 -251.710 -16.430 ;
        RECT -251.490 -17.160 -251.080 -17.040 ;
        RECT -251.990 -17.360 -251.080 -17.160 ;
        RECT -251.990 -17.410 -251.710 -17.360 ;
        RECT -251.970 -17.420 -251.740 -17.410 ;
        RECT -251.490 -17.420 -251.080 -17.360 ;
        RECT -249.020 -17.120 -248.620 -14.870 ;
        RECT -248.120 -17.060 -247.790 -17.000 ;
        RECT -247.500 -17.060 -247.270 -16.400 ;
        RECT -248.120 -17.120 -247.270 -17.060 ;
        RECT -249.020 -17.330 -247.270 -17.120 ;
        RECT -249.020 -17.390 -247.790 -17.330 ;
        RECT -249.020 -17.430 -248.620 -17.390 ;
        RECT -248.120 -17.410 -247.790 -17.390 ;
        RECT -247.500 -17.400 -247.270 -17.330 ;
        RECT -204.530 -37.600 -203.020 -36.910 ;
        RECT -218.160 -37.630 -217.790 -37.600 ;
        RECT -211.640 -37.630 -201.420 -37.600 ;
        RECT -218.160 -37.640 -201.420 -37.630 ;
        RECT -224.720 -37.800 -201.420 -37.640 ;
        RECT -224.720 -44.780 -224.380 -37.800 ;
        RECT -218.160 -37.850 -201.420 -37.800 ;
        RECT -218.160 -38.600 -217.790 -37.850 ;
        RECT -211.640 -37.900 -201.420 -37.850 ;
        RECT -219.160 -38.900 -217.720 -38.600 ;
        RECT -211.630 -39.090 -211.400 -37.900 ;
        RECT -224.780 -44.930 -224.380 -44.780 ;
        RECT -224.720 -44.940 -224.380 -44.930 ;
        RECT -212.310 -39.770 -212.080 -39.710 ;
        RECT -211.670 -39.770 -211.380 -39.090 ;
        RECT -207.530 -39.770 -207.200 -39.060 ;
        RECT -206.800 -39.770 -206.570 -39.660 ;
        RECT -212.310 -40.330 -206.570 -39.770 ;
        RECT -225.810 -46.230 -225.450 -45.220 ;
        RECT -224.720 -47.320 -224.420 -44.940 ;
        RECT -212.310 -47.410 -212.080 -40.330 ;
        RECT -211.670 -40.420 -211.370 -40.330 ;
        RECT -211.630 -40.430 -211.400 -40.420 ;
        RECT -211.680 -47.410 -211.380 -47.330 ;
        RECT -206.800 -47.410 -206.570 -40.330 ;
        RECT -201.720 -40.920 -201.420 -37.900 ;
        RECT -141.330 -38.400 -140.900 27.670 ;
        RECT -99.400 24.530 -97.850 39.150 ;
        RECT -108.930 24.510 -97.850 24.530 ;
        RECT -108.990 23.880 -97.850 24.510 ;
        RECT -108.990 23.840 -108.090 23.880 ;
        RECT -108.990 23.790 -108.680 23.840 ;
        RECT -99.400 21.490 -97.850 23.880 ;
        RECT -39.670 23.230 -37.420 39.150 ;
        RECT 2.330 32.760 3.050 32.820 ;
        RECT 2.310 32.510 3.050 32.760 ;
        RECT 2.310 31.920 3.000 32.510 ;
        RECT 2.310 23.230 2.960 31.920 ;
        RECT -39.910 23.140 5.350 23.230 ;
        RECT 30.450 23.140 31.360 43.310 ;
        RECT 67.150 35.500 67.870 35.810 ;
        RECT 67.230 35.320 67.820 35.500 ;
        RECT 67.180 28.200 67.830 35.320 ;
        RECT 95.580 28.200 96.360 45.850 ;
        RECT 67.180 26.650 96.570 28.200 ;
        RECT 67.180 24.880 67.830 26.650 ;
        RECT 67.000 23.140 67.980 24.880 ;
        RECT -39.910 21.980 68.320 23.140 ;
        RECT -39.910 21.680 5.350 21.980 ;
        RECT -120.380 -3.610 -119.480 -3.055 ;
        RECT -99.310 -3.610 -98.150 21.490 ;
        RECT -39.670 20.720 -35.810 21.680 ;
        RECT -39.640 20.580 -35.810 20.720 ;
        RECT -37.350 12.970 -35.810 20.580 ;
        RECT 10.120 12.970 10.370 12.980 ;
        RECT -37.550 12.280 10.370 12.970 ;
        RECT -120.380 -4.520 -98.150 -3.610 ;
        RECT -120.380 -5.160 -119.480 -4.520 ;
        RECT -159.080 -38.540 -158.770 -38.460 ;
        RECT -159.080 -38.600 -158.180 -38.540 ;
        RECT -141.630 -38.600 -140.840 -38.400 ;
        RECT -159.080 -39.040 -140.840 -38.600 ;
        RECT -159.080 -39.130 -158.180 -39.040 ;
        RECT -159.080 -39.180 -158.770 -39.130 ;
        RECT -141.630 -39.190 -140.840 -39.040 ;
        RECT -99.310 -40.160 -98.150 -4.520 ;
        RECT -111.980 -40.390 -111.670 -40.310 ;
        RECT -101.050 -40.340 -98.150 -40.160 ;
        RECT -111.490 -40.390 -98.150 -40.340 ;
        RECT -111.980 -40.980 -98.150 -40.390 ;
        RECT -111.980 -41.030 -111.670 -40.980 ;
        RECT -111.490 -40.990 -98.150 -40.980 ;
        RECT -212.310 -48.350 -206.570 -47.410 ;
        RECT -212.310 -58.780 -212.080 -48.350 ;
        RECT -211.670 -48.450 -211.380 -48.350 ;
        RECT -211.670 -58.780 -211.370 -58.680 ;
        RECT -206.800 -58.780 -206.570 -48.350 ;
        RECT -212.310 -59.600 -206.570 -58.780 ;
        RECT -212.310 -59.710 -212.080 -59.600 ;
        RECT -211.670 -60.330 -211.380 -59.600 ;
        RECT -206.800 -59.660 -206.570 -59.600 ;
        RECT -122.920 -68.740 -122.020 -67.745 ;
        RECT -104.370 -68.740 -102.820 -40.990 ;
        RECT -101.050 -41.140 -98.150 -40.990 ;
        RECT -99.310 -41.480 -98.150 -41.140 ;
        RECT -37.350 -46.610 -35.810 12.280 ;
        RECT 0.440 4.640 1.040 5.640 ;
        RECT 4.520 4.660 5.120 5.660 ;
        RECT 0.400 1.200 1.000 2.200 ;
        RECT 4.460 1.220 5.060 2.220 ;
        RECT 5.930 -0.470 6.560 -0.300 ;
        RECT 10.120 -0.470 10.370 12.280 ;
        RECT 5.930 -0.620 10.380 -0.470 ;
        RECT 5.930 -0.820 6.560 -0.620 ;
        RECT -37.350 -47.570 -35.000 -46.610 ;
        RECT -37.490 -47.870 7.770 -47.570 ;
        RECT -37.490 -49.030 70.740 -47.870 ;
        RECT -37.490 -49.120 7.770 -49.030 ;
        RECT -122.920 -69.520 -102.820 -68.740 ;
        RECT -122.920 -69.850 -122.020 -69.520 ;
        RECT -104.370 -69.730 -102.820 -69.520 ;
        RECT -37.250 -95.930 -35.000 -49.120 ;
        RECT 4.730 -57.810 5.380 -49.120 ;
        RECT 4.730 -58.400 5.420 -57.810 ;
        RECT 4.730 -58.650 5.470 -58.400 ;
        RECT 4.750 -58.710 5.470 -58.650 ;
        RECT 32.870 -69.200 33.780 -49.030 ;
        RECT 69.420 -50.770 70.400 -49.030 ;
        RECT 69.600 -52.540 70.250 -50.770 ;
        RECT 69.600 -54.090 98.990 -52.540 ;
        RECT 69.600 -61.210 70.250 -54.090 ;
        RECT 69.650 -61.390 70.240 -61.210 ;
        RECT 69.570 -61.700 70.290 -61.390 ;
        RECT 32.315 -70.100 34.420 -69.200 ;
        RECT 98.000 -71.740 98.780 -54.090 ;
        RECT 97.005 -72.640 99.110 -71.740 ;
        RECT 1.150 -90.620 1.590 -89.640 ;
        RECT 67.660 -90.620 68.450 -90.560 ;
        RECT 1.150 -91.050 68.450 -90.620 ;
        RECT 1.150 -93.770 1.590 -91.050 ;
        RECT 67.660 -91.350 68.450 -91.050 ;
        RECT -37.250 -96.030 -21.880 -95.930 ;
        RECT -12.720 -96.030 -7.750 -94.060 ;
        RECT -37.250 -98.410 -7.750 -96.030 ;
        RECT -37.250 -172.610 -35.000 -98.410 ;
        RECT -23.680 -98.510 -7.750 -98.410 ;
        RECT -12.720 -99.720 -7.750 -98.510 ;
        RECT 1.150 -99.490 4.670 -93.770 ;
        RECT 1.150 -106.610 1.590 -99.490 ;
        RECT 1.150 -106.900 1.830 -106.610 ;
        RECT 1.240 -107.200 1.830 -106.900 ;
        RECT 1.160 -107.510 1.880 -107.200 ;
        RECT 67.860 -107.900 68.300 -91.350 ;
        RECT 67.800 -108.490 68.390 -107.900 ;
        RECT 67.720 -108.800 68.440 -108.490 ;
        RECT -32.270 -140.560 -29.460 -135.720 ;
        RECT -31.330 -150.110 -30.490 -140.560 ;
        RECT -31.430 -151.500 -29.050 -150.110 ;
        RECT 66.860 -151.440 70.180 -151.140 ;
        RECT -30.500 -170.510 -29.060 -151.500 ;
        RECT -11.070 -151.870 -7.750 -151.570 ;
        RECT -11.070 -153.440 -10.770 -151.870 ;
        RECT 66.860 -152.740 67.160 -151.440 ;
        RECT -12.390 -155.330 -10.770 -153.440 ;
        RECT 66.170 -154.250 67.160 -152.740 ;
        RECT -11.070 -161.550 -10.770 -155.330 ;
        RECT -9.010 -156.950 10.990 -156.720 ;
        RECT -8.900 -157.350 -8.340 -156.950 ;
        RECT -9.610 -157.680 -8.340 -157.350 ;
        RECT -8.900 -161.520 -8.340 -157.680 ;
        RECT -8.900 -161.530 -8.250 -161.520 ;
        RECT -1.260 -161.530 -0.320 -156.950 ;
        RECT 10.110 -161.520 10.930 -156.950 ;
        RECT 66.860 -161.120 67.160 -154.250 ;
        RECT 68.920 -156.520 88.920 -156.290 ;
        RECT 69.030 -156.920 69.590 -156.520 ;
        RECT 68.320 -157.250 69.590 -156.920 ;
        RECT 69.030 -161.090 69.590 -157.250 ;
        RECT 69.030 -161.100 69.680 -161.090 ;
        RECT 76.670 -161.100 77.610 -156.520 ;
        RECT 88.040 -161.090 88.860 -156.520 ;
        RECT 87.940 -161.100 88.860 -161.090 ;
        RECT 68.350 -161.120 69.680 -161.100 ;
        RECT 66.860 -161.350 69.690 -161.120 ;
        RECT 66.860 -161.360 67.160 -161.350 ;
        RECT 10.010 -161.530 10.930 -161.520 ;
        RECT -9.580 -161.550 -8.250 -161.530 ;
        RECT -11.070 -161.780 -8.240 -161.550 ;
        RECT -11.070 -161.790 -10.770 -161.780 ;
        RECT -11.040 -167.940 -10.820 -161.790 ;
        RECT -9.580 -161.820 -8.250 -161.780 ;
        RECT -1.340 -161.820 -0.220 -161.530 ;
        RECT 10.010 -161.820 11.660 -161.530 ;
        RECT -8.900 -162.230 -8.340 -161.820 ;
        RECT -1.340 -161.830 -0.320 -161.820 ;
        RECT -1.260 -162.230 -0.320 -161.830 ;
        RECT 10.110 -162.230 10.930 -161.820 ;
        RECT -8.960 -162.460 11.040 -162.230 ;
        RECT 66.890 -167.510 67.110 -161.360 ;
        RECT 68.350 -161.390 69.680 -161.350 ;
        RECT 76.590 -161.390 77.710 -161.100 ;
        RECT 87.940 -161.390 89.590 -161.100 ;
        RECT 69.030 -161.800 69.590 -161.390 ;
        RECT 76.590 -161.400 77.610 -161.390 ;
        RECT 76.670 -161.800 77.610 -161.400 ;
        RECT 88.040 -161.800 88.860 -161.390 ;
        RECT 68.970 -162.030 88.970 -161.800 ;
        RECT 67.860 -167.510 68.160 -167.440 ;
        RECT -10.070 -167.940 -9.770 -167.870 ;
        RECT 66.860 -167.880 68.160 -167.510 ;
        RECT -11.070 -168.310 -9.770 -167.940 ;
        RECT -34.750 -172.520 -29.060 -170.510 ;
        RECT -30.500 -205.360 -29.060 -172.520 ;
        RECT -11.030 -174.530 -10.870 -168.310 ;
        RECT -10.070 -169.310 -9.770 -168.310 ;
        RECT 66.900 -174.100 67.060 -167.880 ;
        RECT 67.860 -168.880 68.160 -167.880 ;
        RECT 66.900 -174.140 74.200 -174.100 ;
        RECT 66.900 -174.440 76.580 -174.140 ;
        RECT 74.040 -174.500 74.190 -174.440 ;
        RECT -11.030 -174.570 -3.730 -174.530 ;
        RECT -11.030 -174.870 -1.350 -174.570 ;
        RECT -3.890 -174.930 -3.740 -174.870 ;
        RECT 74.480 -175.530 75.490 -175.170 ;
        RECT -3.450 -175.960 -2.440 -175.600 ;
        RECT 45.660 -197.220 46.660 -196.990 ;
        RECT 46.320 -197.510 46.590 -197.220 ;
        RECT 46.260 -197.840 46.670 -197.510 ;
        RECT 43.670 -198.340 44.130 -198.310 ;
        RECT 46.380 -198.340 46.650 -197.840 ;
        RECT 43.670 -198.740 46.690 -198.340 ;
        RECT 43.670 -201.470 44.130 -198.740 ;
        RECT 46.300 -201.210 46.680 -200.800 ;
        RECT 43.510 -201.500 44.130 -201.470 ;
        RECT 44.680 -201.500 45.050 -201.290 ;
        RECT 46.420 -201.430 46.620 -201.210 ;
        RECT 45.690 -201.460 46.670 -201.430 ;
        RECT 43.510 -202.010 45.050 -201.500 ;
        RECT 45.680 -201.690 46.680 -201.460 ;
        RECT 45.690 -201.710 46.670 -201.690 ;
        RECT 43.510 -203.300 43.830 -202.010 ;
        RECT 44.680 -202.280 45.050 -202.010 ;
        RECT 42.100 -203.810 43.830 -203.300 ;
        RECT 42.100 -204.000 42.650 -203.810 ;
        RECT 39.490 -204.170 42.650 -204.000 ;
        RECT -1.050 -204.270 42.650 -204.170 ;
        RECT -28.800 -204.940 42.650 -204.270 ;
        RECT -28.800 -205.020 39.750 -204.940 ;
        RECT -28.800 -205.120 12.000 -205.020 ;
        RECT 42.100 -223.590 42.650 -204.940 ;
        RECT 43.510 -205.030 43.830 -203.810 ;
        RECT 44.860 -204.840 45.170 -204.800 ;
        RECT 44.850 -205.030 45.170 -204.840 ;
        RECT 43.510 -205.610 45.170 -205.030 ;
        RECT 43.510 -205.650 43.830 -205.610 ;
        RECT 44.850 -205.700 45.170 -205.610 ;
        RECT 44.860 -205.740 45.170 -205.700 ;
        RECT 45.500 -217.510 46.500 -217.280 ;
        RECT 46.160 -217.800 46.430 -217.510 ;
        RECT 46.100 -218.130 46.510 -217.800 ;
        RECT 43.510 -218.630 43.970 -218.600 ;
        RECT 46.220 -218.630 46.490 -218.130 ;
        RECT 43.510 -219.030 46.530 -218.630 ;
        RECT 43.510 -221.760 43.970 -219.030 ;
        RECT 46.140 -221.500 46.520 -221.090 ;
        RECT 43.350 -221.790 43.970 -221.760 ;
        RECT 44.520 -221.790 44.890 -221.580 ;
        RECT 46.260 -221.720 46.460 -221.500 ;
        RECT 45.530 -221.750 46.510 -221.720 ;
        RECT 43.350 -222.300 44.890 -221.790 ;
        RECT 45.520 -221.980 46.520 -221.750 ;
        RECT 45.530 -222.000 46.510 -221.980 ;
        RECT 43.350 -223.590 43.670 -222.300 ;
        RECT 44.520 -222.570 44.890 -222.300 ;
        RECT 42.010 -224.100 43.670 -223.590 ;
        RECT 42.100 -224.210 42.690 -224.100 ;
        RECT 42.410 -237.520 42.690 -224.210 ;
        RECT 43.350 -225.320 43.670 -224.100 ;
        RECT 44.700 -225.130 45.010 -225.090 ;
        RECT 44.690 -225.320 45.010 -225.130 ;
        RECT 43.350 -225.900 45.010 -225.320 ;
        RECT 43.350 -225.940 43.670 -225.900 ;
        RECT 44.690 -225.990 45.010 -225.900 ;
        RECT 44.700 -226.030 45.010 -225.990 ;
        RECT 44.600 -237.270 45.600 -237.040 ;
        RECT 45.270 -237.520 45.520 -237.270 ;
        RECT 42.410 -237.570 45.570 -237.520 ;
        RECT 42.410 -237.900 45.610 -237.570 ;
      LAYER via ;
        RECT -98.570 71.010 -97.350 72.040 ;
        RECT -14.250 128.310 -13.950 128.900 ;
        RECT 64.040 127.570 64.300 127.930 ;
        RECT -33.550 112.050 -33.020 112.670 ;
        RECT -13.390 70.400 -11.820 72.490 ;
        RECT -188.840 59.860 -188.220 60.390 ;
        RECT -205.070 40.790 -204.480 41.090 ;
        RECT -148.660 38.660 -146.570 40.230 ;
        RECT -0.220 70.350 0.760 71.980 ;
        RECT -148.150 26.080 -146.520 27.060 ;
        RECT -204.100 -37.460 -203.740 -37.200 ;
        RECT 0.540 4.740 0.940 5.540 ;
        RECT 4.620 4.760 5.020 5.560 ;
        RECT 0.500 1.300 0.900 2.100 ;
        RECT 4.560 1.320 4.960 2.120 ;
        RECT 6.120 -0.640 6.380 -0.380 ;
        RECT -10.970 -98.380 -9.400 -96.290 ;
        RECT 2.200 -97.870 3.180 -96.240 ;
        RECT -31.130 -138.560 -30.600 -137.940 ;
        RECT -11.830 -154.790 -11.530 -154.200 ;
        RECT 66.460 -153.820 66.720 -153.460 ;
      LAYER met2 ;
        RECT -365.150 -323.900 -355.150 301.100 ;
        RECT -99.100 72.860 -96.770 301.060 ;
        RECT -14.540 127.830 -13.630 129.280 ;
        RECT 63.040 127.980 63.310 128.010 ;
        RECT 63.860 127.980 64.430 128.240 ;
        RECT -14.340 121.180 -13.860 127.830 ;
        RECT 63.040 127.580 64.430 127.980 ;
        RECT -14.490 113.090 -13.740 121.180 ;
        RECT -34.390 111.490 -13.740 113.090 ;
        RECT -14.490 108.900 -13.740 111.490 ;
        RECT -14.490 108.880 62.790 108.900 ;
        RECT 63.040 108.880 63.310 127.580 ;
        RECT 63.860 126.990 64.430 127.580 ;
        RECT -14.490 108.230 63.350 108.880 ;
        RECT -14.060 108.190 63.350 108.230 ;
        RECT 62.720 108.160 63.350 108.190 ;
        RECT -99.670 70.150 -96.060 72.860 ;
        RECT -14.780 72.280 -10.650 73.230 ;
        RECT -1.000 72.280 1.860 73.170 ;
        RECT -14.780 70.180 1.860 72.280 ;
        RECT -14.780 68.700 -10.650 70.180 ;
        RECT -1.000 68.230 1.860 70.180 ;
        RECT -205.450 41.180 -204.000 41.380 ;
        RECT -189.260 41.330 -187.660 61.230 ;
        RECT -197.350 41.180 -184.400 41.330 ;
        RECT -205.450 40.900 -184.400 41.180 ;
        RECT -205.450 40.700 -184.360 40.900 ;
        RECT -205.450 40.470 -204.000 40.700 ;
        RECT -197.350 40.580 -184.360 40.700 ;
        RECT -185.070 -35.880 -184.360 40.580 ;
        RECT -149.400 37.490 -144.870 41.620 ;
        RECT -148.450 27.840 -146.350 37.490 ;
        RECT -149.340 24.980 -144.400 27.840 ;
        RECT 0.440 3.840 1.040 6.240 ;
        RECT 4.515 3.860 5.120 6.260 ;
        RECT 0.440 2.800 1.000 3.840 ;
        RECT 4.515 2.820 5.060 3.860 ;
        RECT 0.400 0.400 1.000 2.800 ;
        RECT 4.460 0.420 5.060 2.820 ;
        RECT 0.520 -0.460 0.910 0.400 ;
        RECT 4.550 -0.460 4.940 0.420 ;
        RECT 5.960 -0.460 6.530 -0.330 ;
        RECT 0.520 -0.660 6.530 -0.460 ;
        RECT 0.530 -0.670 6.530 -0.660 ;
        RECT 5.960 -0.780 6.530 -0.670 ;
        RECT -185.070 -35.950 -184.330 -35.880 ;
        RECT -185.050 -36.200 -184.330 -35.950 ;
        RECT -204.180 -36.470 -184.330 -36.200 ;
        RECT -204.150 -37.020 -203.750 -36.470 ;
        RECT -185.050 -36.510 -184.330 -36.470 ;
        RECT -204.410 -37.590 -203.160 -37.020 ;
        RECT -12.360 -96.070 -8.230 -94.590 ;
        RECT 1.420 -96.070 4.280 -94.120 ;
        RECT -12.360 -98.170 4.280 -96.070 ;
        RECT -12.360 -99.120 -8.230 -98.170 ;
        RECT 1.420 -99.060 4.280 -98.170 ;
        RECT 65.140 -134.080 65.770 -134.050 ;
        RECT -11.640 -134.120 65.770 -134.080 ;
        RECT -12.070 -134.770 65.770 -134.120 ;
        RECT -12.070 -134.790 65.210 -134.770 ;
        RECT -12.070 -137.380 -11.320 -134.790 ;
        RECT -31.970 -138.980 -11.320 -137.380 ;
        RECT -12.070 -147.070 -11.320 -138.980 ;
        RECT -11.920 -153.720 -11.440 -147.070 ;
        RECT 65.460 -153.470 65.730 -134.770 ;
        RECT 66.280 -153.470 66.850 -152.880 ;
        RECT -12.120 -155.170 -11.210 -153.720 ;
        RECT 65.460 -153.870 66.850 -153.470 ;
        RECT 65.460 -153.900 65.730 -153.870 ;
        RECT 66.280 -154.130 66.850 -153.870 ;
        RECT 204.850 -323.900 214.850 301.100 ;
      LAYER via2 ;
        RECT -362.650 293.600 -357.650 298.600 ;
        RECT -98.520 292.050 -97.230 300.370 ;
        RECT 207.350 293.600 212.350 298.600 ;
        RECT -362.650 -321.400 -357.650 -316.400 ;
        RECT 207.350 -321.400 212.350 -316.400 ;
      LAYER met3 ;
        RECT -400.150 291.100 249.850 301.100 ;
        RECT -400.150 -323.900 249.850 -313.900 ;
    END
  END vssd1
  PIN vccd1
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 44.450 209.940 47.640 212.050 ;
        RECT 45.800 198.580 48.990 200.690 ;
        RECT 45.820 195.160 49.010 197.270 ;
        RECT 45.890 190.170 49.080 192.280 ;
        RECT 45.960 178.290 49.150 180.400 ;
        RECT 45.980 174.870 49.170 176.980 ;
        RECT 46.050 169.880 49.240 171.990 ;
        RECT -2.610 148.530 0.580 150.640 ;
        RECT 75.320 148.100 78.510 150.210 ;
        RECT -226.810 26.260 -224.700 29.450 ;
        RECT -288.220 -20.800 -286.110 -17.610 ;
        RECT -276.860 -22.150 -274.750 -18.960 ;
        RECT -273.440 -22.170 -271.330 -18.980 ;
        RECT -268.450 -22.240 -266.340 -19.050 ;
        RECT -256.570 -22.310 -254.460 -19.120 ;
        RECT -253.150 -22.330 -251.040 -19.140 ;
        RECT -248.160 -22.400 -246.050 -19.210 ;
        RECT -226.380 -51.670 -224.270 -48.480 ;
        RECT -0.190 -176.530 3.000 -174.420 ;
        RECT 77.740 -176.100 80.930 -173.990 ;
        RECT 48.470 -197.880 51.660 -195.770 ;
        RECT 48.400 -202.870 51.590 -200.760 ;
        RECT 48.380 -206.290 51.570 -204.180 ;
        RECT 48.310 -218.170 51.500 -216.060 ;
        RECT 48.240 -223.160 51.430 -221.050 ;
        RECT 48.220 -226.580 51.410 -224.470 ;
        RECT 46.870 -237.940 50.060 -235.830 ;
      LAYER li1 ;
        RECT 44.630 211.700 47.460 211.870 ;
        RECT 44.630 210.290 44.800 211.700 ;
        RECT 45.525 211.130 46.565 211.300 ;
        RECT 47.290 210.290 47.460 211.700 ;
        RECT 44.630 210.120 47.460 210.290 ;
        RECT 45.980 200.340 48.810 200.510 ;
        RECT 45.980 198.930 46.150 200.340 ;
        RECT 46.875 199.330 47.915 199.500 ;
        RECT 48.640 198.930 48.810 200.340 ;
        RECT 45.980 198.760 48.810 198.930 ;
        RECT 46.000 196.920 48.830 197.090 ;
        RECT 46.000 195.510 46.170 196.920 ;
        RECT 46.895 196.350 47.935 196.520 ;
        RECT 48.660 195.510 48.830 196.920 ;
        RECT 46.000 195.340 48.830 195.510 ;
        RECT 46.070 191.930 48.900 192.100 ;
        RECT 46.070 190.520 46.240 191.930 ;
        RECT 46.965 191.360 48.005 191.530 ;
        RECT 48.730 190.520 48.900 191.930 ;
        RECT 46.070 190.350 48.900 190.520 ;
        RECT 46.140 180.050 48.970 180.220 ;
        RECT 46.140 178.640 46.310 180.050 ;
        RECT 47.035 179.040 48.075 179.210 ;
        RECT 48.800 178.640 48.970 180.050 ;
        RECT 46.140 178.470 48.970 178.640 ;
        RECT 46.160 176.630 48.990 176.800 ;
        RECT 46.160 175.220 46.330 176.630 ;
        RECT 47.055 176.060 48.095 176.230 ;
        RECT 48.820 175.220 48.990 176.630 ;
        RECT 46.160 175.050 48.990 175.220 ;
        RECT 46.230 171.640 49.060 171.810 ;
        RECT 46.230 170.230 46.400 171.640 ;
        RECT 47.125 171.070 48.165 171.240 ;
        RECT 48.890 170.230 49.060 171.640 ;
        RECT 46.230 170.060 49.060 170.230 ;
        RECT -2.430 150.290 0.400 150.460 ;
        RECT -2.430 148.880 -2.260 150.290 ;
        RECT -1.460 149.890 -0.570 150.290 ;
        RECT -1.535 149.720 -0.495 149.890 ;
        RECT 0.230 148.880 0.400 150.290 ;
        RECT -2.430 148.710 0.400 148.880 ;
        RECT 75.500 149.860 78.330 150.030 ;
        RECT 75.500 148.450 75.670 149.860 ;
        RECT 76.470 149.460 77.360 149.860 ;
        RECT 76.395 149.290 77.435 149.460 ;
        RECT 78.160 148.450 78.330 149.860 ;
        RECT 75.500 148.280 78.330 148.450 ;
        RECT -226.630 29.100 -224.880 29.270 ;
        RECT -226.630 28.300 -226.460 29.100 ;
        RECT -226.060 28.300 -225.890 28.375 ;
        RECT -226.630 27.410 -225.890 28.300 ;
        RECT -226.630 26.610 -226.460 27.410 ;
        RECT -226.060 27.335 -225.890 27.410 ;
        RECT -225.050 26.610 -224.880 29.100 ;
        RECT -226.630 26.440 -224.880 26.610 ;
        RECT -288.040 -17.960 -286.290 -17.790 ;
        RECT -288.040 -20.450 -287.870 -17.960 ;
        RECT -287.470 -19.725 -287.300 -18.685 ;
        RECT -286.460 -20.450 -286.290 -17.960 ;
        RECT -288.040 -20.620 -286.290 -20.450 ;
        RECT -276.680 -19.310 -274.930 -19.140 ;
        RECT -276.680 -21.800 -276.510 -19.310 ;
        RECT -275.670 -21.075 -275.500 -20.035 ;
        RECT -275.100 -21.800 -274.930 -19.310 ;
        RECT -276.680 -21.970 -274.930 -21.800 ;
        RECT -273.260 -19.330 -271.510 -19.160 ;
        RECT -273.260 -21.820 -273.090 -19.330 ;
        RECT -272.690 -21.095 -272.520 -20.055 ;
        RECT -271.680 -21.820 -271.510 -19.330 ;
        RECT -273.260 -21.990 -271.510 -21.820 ;
        RECT -268.270 -19.400 -266.520 -19.230 ;
        RECT -268.270 -21.890 -268.100 -19.400 ;
        RECT -267.700 -21.165 -267.530 -20.125 ;
        RECT -266.690 -21.890 -266.520 -19.400 ;
        RECT -268.270 -22.060 -266.520 -21.890 ;
        RECT -256.390 -19.470 -254.640 -19.300 ;
        RECT -256.390 -21.960 -256.220 -19.470 ;
        RECT -255.380 -21.235 -255.210 -20.195 ;
        RECT -254.810 -21.960 -254.640 -19.470 ;
        RECT -256.390 -22.130 -254.640 -21.960 ;
        RECT -252.970 -19.490 -251.220 -19.320 ;
        RECT -252.970 -21.980 -252.800 -19.490 ;
        RECT -252.400 -21.255 -252.230 -20.215 ;
        RECT -251.390 -21.980 -251.220 -19.490 ;
        RECT -252.970 -22.150 -251.220 -21.980 ;
        RECT -247.980 -19.560 -246.230 -19.390 ;
        RECT -247.980 -22.050 -247.810 -19.560 ;
        RECT -247.410 -21.325 -247.240 -20.285 ;
        RECT -246.400 -22.050 -246.230 -19.560 ;
        RECT -247.980 -22.220 -246.230 -22.050 ;
        RECT -226.200 -48.830 -224.450 -48.660 ;
        RECT -226.200 -49.630 -226.030 -48.830 ;
        RECT -225.630 -49.630 -225.460 -49.555 ;
        RECT -226.200 -50.520 -225.460 -49.630 ;
        RECT -226.200 -51.320 -226.030 -50.520 ;
        RECT -225.630 -50.595 -225.460 -50.520 ;
        RECT -224.620 -51.320 -224.450 -48.830 ;
        RECT -226.200 -51.490 -224.450 -51.320 ;
        RECT 77.920 -174.340 80.750 -174.170 ;
        RECT -0.010 -174.770 2.820 -174.600 ;
        RECT -0.010 -176.180 0.160 -174.770 ;
        RECT 0.885 -175.780 1.925 -175.610 ;
        RECT 0.960 -176.180 1.850 -175.780 ;
        RECT 2.650 -176.180 2.820 -174.770 ;
        RECT 77.920 -175.750 78.090 -174.340 ;
        RECT 78.815 -175.350 79.855 -175.180 ;
        RECT 78.890 -175.750 79.780 -175.350 ;
        RECT 80.580 -175.750 80.750 -174.340 ;
        RECT 77.920 -175.920 80.750 -175.750 ;
        RECT -0.010 -176.350 2.820 -176.180 ;
        RECT 48.650 -196.120 51.480 -195.950 ;
        RECT 48.650 -197.530 48.820 -196.120 ;
        RECT 49.545 -197.130 50.585 -196.960 ;
        RECT 51.310 -197.530 51.480 -196.120 ;
        RECT 48.650 -197.700 51.480 -197.530 ;
        RECT 48.580 -201.110 51.410 -200.940 ;
        RECT 48.580 -202.520 48.750 -201.110 ;
        RECT 49.475 -202.120 50.515 -201.950 ;
        RECT 51.240 -202.520 51.410 -201.110 ;
        RECT 48.580 -202.690 51.410 -202.520 ;
        RECT 48.560 -204.530 51.390 -204.360 ;
        RECT 48.560 -205.940 48.730 -204.530 ;
        RECT 49.455 -205.100 50.495 -204.930 ;
        RECT 51.220 -205.940 51.390 -204.530 ;
        RECT 48.560 -206.110 51.390 -205.940 ;
        RECT 48.490 -216.410 51.320 -216.240 ;
        RECT 48.490 -217.820 48.660 -216.410 ;
        RECT 49.385 -217.420 50.425 -217.250 ;
        RECT 51.150 -217.820 51.320 -216.410 ;
        RECT 48.490 -217.990 51.320 -217.820 ;
        RECT 48.420 -221.400 51.250 -221.230 ;
        RECT 48.420 -222.810 48.590 -221.400 ;
        RECT 49.315 -222.410 50.355 -222.240 ;
        RECT 51.080 -222.810 51.250 -221.400 ;
        RECT 48.420 -222.980 51.250 -222.810 ;
        RECT 48.400 -224.820 51.230 -224.650 ;
        RECT 48.400 -226.230 48.570 -224.820 ;
        RECT 49.295 -225.390 50.335 -225.220 ;
        RECT 51.060 -226.230 51.230 -224.820 ;
        RECT 48.400 -226.400 51.230 -226.230 ;
        RECT 47.050 -236.180 49.880 -236.010 ;
        RECT 47.050 -237.590 47.220 -236.180 ;
        RECT 47.945 -237.190 48.985 -237.020 ;
        RECT 49.710 -237.590 49.880 -236.180 ;
        RECT 47.050 -237.760 49.880 -237.590 ;
      LAYER mcon ;
        RECT 46.060 211.700 46.490 211.870 ;
        RECT 45.605 211.130 46.485 211.300 ;
        RECT 46.955 199.330 47.835 199.500 ;
        RECT 47.430 198.760 47.830 198.930 ;
        RECT 47.510 196.920 47.810 197.090 ;
        RECT 46.975 196.350 47.855 196.520 ;
        RECT 47.690 191.930 47.930 192.100 ;
        RECT 47.045 191.360 47.925 191.530 ;
        RECT 47.115 179.040 47.995 179.210 ;
        RECT 47.590 178.470 47.990 178.640 ;
        RECT 47.670 176.630 47.970 176.800 ;
        RECT 47.135 176.060 48.015 176.230 ;
        RECT 47.850 171.640 48.090 171.810 ;
        RECT 47.205 171.070 48.085 171.240 ;
        RECT -1.455 149.720 -0.575 149.890 ;
        RECT -1.950 148.710 -0.080 148.880 ;
        RECT 76.475 149.290 77.355 149.460 ;
        RECT 75.980 148.280 77.850 148.450 ;
        RECT -226.060 27.415 -225.890 28.295 ;
        RECT -225.050 26.920 -224.880 28.790 ;
        RECT -288.040 -19.650 -287.870 -19.220 ;
        RECT -287.470 -19.645 -287.300 -18.765 ;
        RECT -275.670 -20.995 -275.500 -20.115 ;
        RECT -275.100 -20.990 -274.930 -20.590 ;
        RECT -273.260 -20.970 -273.090 -20.670 ;
        RECT -272.690 -21.015 -272.520 -20.135 ;
        RECT -268.270 -21.090 -268.100 -20.850 ;
        RECT -267.700 -21.085 -267.530 -20.205 ;
        RECT -255.380 -21.155 -255.210 -20.275 ;
        RECT -254.810 -21.150 -254.640 -20.750 ;
        RECT -252.970 -21.130 -252.800 -20.830 ;
        RECT -252.400 -21.175 -252.230 -20.295 ;
        RECT -247.980 -21.250 -247.810 -21.010 ;
        RECT -247.410 -21.245 -247.240 -20.365 ;
        RECT -225.630 -50.515 -225.460 -49.635 ;
        RECT -224.620 -51.010 -224.450 -49.140 ;
        RECT 78.400 -174.340 80.270 -174.170 ;
        RECT 0.470 -174.770 2.340 -174.600 ;
        RECT 0.965 -175.780 1.845 -175.610 ;
        RECT 78.895 -175.350 79.775 -175.180 ;
        RECT 49.625 -197.130 50.505 -196.960 ;
        RECT 50.270 -197.700 50.510 -197.530 ;
        RECT 49.555 -202.120 50.435 -201.950 ;
        RECT 50.090 -202.690 50.390 -202.520 ;
        RECT 50.010 -204.530 50.410 -204.360 ;
        RECT 49.535 -205.100 50.415 -204.930 ;
        RECT 49.465 -217.420 50.345 -217.250 ;
        RECT 50.110 -217.990 50.350 -217.820 ;
        RECT 49.395 -222.410 50.275 -222.240 ;
        RECT 49.930 -222.980 50.230 -222.810 ;
        RECT 49.850 -224.820 50.250 -224.650 ;
        RECT 49.375 -225.390 50.255 -225.220 ;
        RECT 48.025 -237.190 48.905 -237.020 ;
        RECT 48.480 -237.760 48.910 -237.590 ;
      LAYER met1 ;
        RECT 52.100 211.970 52.790 212.080 ;
        RECT 46.060 211.950 52.790 211.970 ;
        RECT 45.960 211.650 52.790 211.950 ;
        RECT 46.060 211.570 52.790 211.650 ;
        RECT 46.070 211.330 46.490 211.570 ;
        RECT 45.545 211.100 46.545 211.330 ;
        RECT 46.895 199.300 47.895 199.530 ;
        RECT 47.430 199.010 47.830 199.300 ;
        RECT 47.370 198.660 47.890 199.010 ;
        RECT 47.540 198.140 47.810 198.660 ;
        RECT 49.420 198.190 50.620 198.200 ;
        RECT 49.420 198.140 50.640 198.190 ;
        RECT 47.540 197.760 50.640 198.140 ;
        RECT 47.540 197.150 47.810 197.760 ;
        RECT 49.420 197.720 50.640 197.760 ;
        RECT 47.440 196.870 47.880 197.150 ;
        RECT 47.490 196.550 47.810 196.870 ;
        RECT 46.915 196.320 47.915 196.550 ;
        RECT 50.440 196.420 50.640 197.720 ;
        RECT 52.100 196.450 52.790 211.570 ;
        RECT 57.710 196.550 58.410 196.570 ;
        RECT 53.690 196.450 58.410 196.550 ;
        RECT 51.330 196.420 58.410 196.450 ;
        RECT 50.440 195.670 58.410 196.420 ;
        RECT 50.440 192.920 50.640 195.670 ;
        RECT 51.330 195.660 58.410 195.670 ;
        RECT 51.330 195.610 53.700 195.660 ;
        RECT 52.100 195.480 52.790 195.610 ;
        RECT 47.660 192.470 50.740 192.920 ;
        RECT 47.680 192.180 47.930 192.470 ;
        RECT 47.600 191.810 48.010 192.180 ;
        RECT 47.680 191.560 47.930 191.810 ;
        RECT 46.985 191.330 47.985 191.560 ;
        RECT 57.710 190.750 58.410 195.660 ;
        RECT 85.960 190.920 86.280 191.070 ;
        RECT 59.790 190.750 86.320 190.920 ;
        RECT 57.710 189.910 86.320 190.750 ;
        RECT 57.710 189.860 60.530 189.910 ;
        RECT 47.055 179.010 48.055 179.240 ;
        RECT 47.590 178.720 47.990 179.010 ;
        RECT 47.530 178.370 48.050 178.720 ;
        RECT 47.700 177.850 47.970 178.370 ;
        RECT 49.580 177.900 50.780 177.910 ;
        RECT 49.580 177.850 50.800 177.900 ;
        RECT 47.700 177.470 50.800 177.850 ;
        RECT 47.700 176.860 47.970 177.470 ;
        RECT 49.580 177.430 50.800 177.470 ;
        RECT 47.600 176.580 48.040 176.860 ;
        RECT 47.650 176.260 47.970 176.580 ;
        RECT 47.075 176.030 48.075 176.260 ;
        RECT 50.600 176.130 50.800 177.430 ;
        RECT 57.710 176.170 58.410 189.860 ;
        RECT 56.130 176.150 58.410 176.170 ;
        RECT 51.750 176.130 58.410 176.150 ;
        RECT 50.600 175.380 58.410 176.130 ;
        RECT 50.600 172.630 50.800 175.380 ;
        RECT 51.750 175.370 58.410 175.380 ;
        RECT 56.130 175.280 58.410 175.370 ;
        RECT 57.710 175.150 58.410 175.280 ;
        RECT 85.960 176.950 86.280 189.910 ;
        RECT 89.260 176.950 90.410 177.320 ;
        RECT 85.960 176.660 90.410 176.950 ;
        RECT 47.820 172.180 50.900 172.630 ;
        RECT 47.840 171.890 48.090 172.180 ;
        RECT 47.760 171.520 48.170 171.890 ;
        RECT 47.840 171.270 48.090 171.520 ;
        RECT 47.145 171.040 48.145 171.270 ;
        RECT 82.330 166.850 84.620 167.920 ;
        RECT 85.960 166.870 86.280 176.660 ;
        RECT 89.260 176.110 90.410 176.660 ;
        RECT 85.760 166.850 86.280 166.870 ;
        RECT 82.330 166.010 86.280 166.850 ;
        RECT 82.330 164.170 84.620 166.010 ;
        RECT 85.150 165.730 86.280 166.010 ;
        RECT 50.670 155.860 51.980 157.300 ;
        RECT -1.510 149.920 -0.520 150.030 ;
        RECT -1.515 149.690 -0.515 149.920 ;
        RECT -1.510 149.680 -0.520 149.690 ;
        RECT -1.500 149.660 -0.520 149.680 ;
        RECT -2.660 148.920 0.030 148.980 ;
        RECT -2.660 148.890 0.550 148.920 ;
        RECT 51.260 148.890 51.750 155.860 ;
        RECT 76.420 149.490 77.410 149.600 ;
        RECT 76.415 149.260 77.415 149.490 ;
        RECT 76.420 149.250 77.410 149.260 ;
        RECT 76.430 149.230 77.410 149.250 ;
        RECT -2.660 148.740 51.750 148.890 ;
        RECT -2.660 148.700 0.550 148.740 ;
        RECT -2.660 148.680 0.030 148.700 ;
        RECT 51.260 148.620 51.750 148.740 ;
        RECT 75.270 148.490 77.960 148.550 ;
        RECT 75.270 148.460 82.000 148.490 ;
        RECT 85.150 148.460 85.750 165.730 ;
        RECT 75.270 148.250 85.750 148.460 ;
        RECT 77.560 148.240 85.750 148.250 ;
        RECT 80.950 148.210 85.750 148.240 ;
        RECT 85.150 148.090 85.750 148.210 ;
        RECT -226.090 28.350 -225.860 28.355 ;
        RECT -226.200 28.340 -225.850 28.350 ;
        RECT -226.200 27.360 -225.830 28.340 ;
        RECT -226.090 27.355 -225.860 27.360 ;
        RECT -225.150 26.810 -224.850 29.500 ;
        RECT -225.090 26.290 -224.870 26.810 ;
        RECT -288.120 -19.220 -287.820 -19.120 ;
        RECT -288.140 -19.230 -287.740 -19.220 ;
        RECT -287.500 -19.230 -287.270 -18.705 ;
        RECT -288.140 -19.650 -287.270 -19.230 ;
        RECT -288.140 -25.260 -287.740 -19.650 ;
        RECT -287.500 -19.705 -287.270 -19.650 ;
        RECT -275.700 -20.590 -275.470 -20.055 ;
        RECT -275.180 -20.590 -274.830 -20.530 ;
        RECT -275.700 -20.700 -274.830 -20.590 ;
        RECT -273.320 -20.650 -273.040 -20.600 ;
        RECT -272.720 -20.650 -272.490 -20.075 ;
        RECT -273.320 -20.700 -272.490 -20.650 ;
        RECT -275.700 -20.970 -272.490 -20.700 ;
        RECT -275.700 -20.990 -274.830 -20.970 ;
        RECT -275.700 -21.055 -275.470 -20.990 ;
        RECT -275.180 -21.050 -274.830 -20.990 ;
        RECT -274.310 -22.580 -273.930 -20.970 ;
        RECT -273.320 -21.040 -273.040 -20.970 ;
        RECT -272.720 -21.075 -272.490 -20.970 ;
        RECT -269.090 -20.840 -268.640 -20.820 ;
        RECT -268.350 -20.840 -267.980 -20.760 ;
        RECT -267.730 -20.840 -267.500 -20.145 ;
        RECT -269.090 -21.090 -267.500 -20.840 ;
        RECT -274.370 -23.600 -273.890 -22.580 ;
        RECT -269.090 -23.600 -268.640 -21.090 ;
        RECT -268.350 -21.170 -267.980 -21.090 ;
        RECT -267.730 -21.145 -267.500 -21.090 ;
        RECT -255.410 -20.750 -255.180 -20.215 ;
        RECT -254.890 -20.750 -254.540 -20.690 ;
        RECT -255.410 -20.860 -254.540 -20.750 ;
        RECT -253.030 -20.810 -252.750 -20.760 ;
        RECT -252.430 -20.810 -252.200 -20.235 ;
        RECT -253.030 -20.860 -252.200 -20.810 ;
        RECT -255.410 -21.130 -252.200 -20.860 ;
        RECT -255.410 -21.150 -254.540 -21.130 ;
        RECT -255.410 -21.215 -255.180 -21.150 ;
        RECT -254.890 -21.210 -254.540 -21.150 ;
        RECT -254.020 -22.740 -253.640 -21.130 ;
        RECT -253.030 -21.200 -252.750 -21.130 ;
        RECT -252.430 -21.235 -252.200 -21.130 ;
        RECT -248.800 -21.000 -248.350 -20.980 ;
        RECT -248.060 -21.000 -247.690 -20.920 ;
        RECT -247.440 -21.000 -247.210 -20.305 ;
        RECT -248.800 -21.250 -247.210 -21.000 ;
        RECT -274.370 -23.780 -268.640 -23.600 ;
        RECT -274.360 -23.800 -268.640 -23.780 ;
        RECT -272.590 -24.490 -271.840 -23.800 ;
        RECT -269.090 -23.900 -268.640 -23.800 ;
        RECT -254.080 -23.760 -253.600 -22.740 ;
        RECT -248.800 -23.760 -248.350 -21.250 ;
        RECT -248.060 -21.330 -247.690 -21.250 ;
        RECT -247.440 -21.305 -247.210 -21.250 ;
        RECT -254.080 -23.940 -248.350 -23.760 ;
        RECT -254.070 -23.960 -248.350 -23.940 ;
        RECT -272.620 -25.260 -271.780 -24.490 ;
        RECT -252.300 -24.910 -251.550 -23.960 ;
        RECT -248.800 -24.060 -248.350 -23.960 ;
        RECT -233.470 -24.420 -232.030 -23.830 ;
        RECT -225.060 -24.420 -224.910 26.290 ;
        RECT -233.470 -24.910 -224.790 -24.420 ;
        RECT -288.250 -25.950 -271.650 -25.260 ;
        RECT -272.620 -26.850 -271.780 -25.950 ;
        RECT -272.720 -26.860 -271.780 -26.850 ;
        RECT -272.720 -30.870 -271.830 -26.860 ;
        RECT -252.320 -29.290 -251.540 -24.910 ;
        RECT -233.470 -25.140 -232.030 -24.910 ;
        RECT -252.340 -30.870 -251.450 -29.290 ;
        RECT -272.740 -31.570 -251.320 -30.870 ;
        RECT -266.920 -32.950 -266.030 -31.570 ;
        RECT -267.090 -33.690 -266.030 -32.950 ;
        RECT -267.090 -59.120 -266.080 -33.690 ;
        RECT -225.660 -49.580 -225.430 -49.575 ;
        RECT -225.770 -49.590 -225.420 -49.580 ;
        RECT -225.770 -50.570 -225.400 -49.590 ;
        RECT -225.660 -50.575 -225.430 -50.570 ;
        RECT -224.720 -50.720 -224.420 -48.430 ;
        RECT -224.720 -51.120 -224.410 -50.720 ;
        RECT -224.660 -54.110 -224.410 -51.120 ;
        RECT -224.660 -55.160 -224.380 -54.110 ;
        RECT -244.090 -57.780 -240.340 -55.490 ;
        RECT -243.020 -58.310 -242.180 -57.780 ;
        RECT -224.630 -58.310 -224.380 -55.160 ;
        RECT -243.020 -58.910 -224.260 -58.310 ;
        RECT -243.020 -58.920 -241.900 -58.910 ;
        RECT -243.040 -59.120 -241.900 -58.920 ;
        RECT -267.240 -59.440 -241.900 -59.120 ;
        RECT -267.090 -59.480 -266.080 -59.440 ;
        RECT -253.120 -62.360 -252.830 -59.440 ;
        RECT -253.240 -62.810 -252.690 -62.360 ;
        RECT 87.570 -174.100 88.170 -173.980 ;
        RECT 83.370 -174.130 88.170 -174.100 ;
        RECT 79.980 -174.140 88.170 -174.130 ;
        RECT 77.690 -174.350 88.170 -174.140 ;
        RECT 77.690 -174.380 84.420 -174.350 ;
        RECT 77.690 -174.440 80.380 -174.380 ;
        RECT -0.240 -174.590 2.450 -174.570 ;
        RECT -0.240 -174.630 2.970 -174.590 ;
        RECT 53.680 -174.630 54.170 -174.510 ;
        RECT -0.240 -174.780 54.170 -174.630 ;
        RECT -0.240 -174.810 2.970 -174.780 ;
        RECT -0.240 -174.870 2.450 -174.810 ;
        RECT 0.920 -175.570 1.900 -175.550 ;
        RECT 0.910 -175.580 1.900 -175.570 ;
        RECT 0.905 -175.810 1.905 -175.580 ;
        RECT 0.910 -175.920 1.900 -175.810 ;
        RECT 53.680 -181.750 54.170 -174.780 ;
        RECT 78.850 -175.140 79.830 -175.120 ;
        RECT 78.840 -175.150 79.830 -175.140 ;
        RECT 78.835 -175.380 79.835 -175.150 ;
        RECT 78.840 -175.490 79.830 -175.380 ;
        RECT 53.090 -183.190 54.400 -181.750 ;
        RECT 84.750 -191.900 87.040 -190.060 ;
        RECT 87.570 -191.620 88.170 -174.350 ;
        RECT 87.570 -191.900 88.700 -191.620 ;
        RECT 84.750 -192.740 88.700 -191.900 ;
        RECT 84.750 -193.810 87.040 -192.740 ;
        RECT 88.180 -192.760 88.700 -192.740 ;
        RECT 49.565 -197.160 50.565 -196.930 ;
        RECT 50.260 -197.410 50.510 -197.160 ;
        RECT 50.180 -197.780 50.590 -197.410 ;
        RECT 50.260 -198.070 50.510 -197.780 ;
        RECT 50.240 -198.520 53.320 -198.070 ;
        RECT 53.020 -201.270 53.220 -198.520 ;
        RECT 60.130 -201.170 60.830 -201.040 ;
        RECT 58.550 -201.260 60.830 -201.170 ;
        RECT 54.170 -201.270 60.830 -201.260 ;
        RECT 49.495 -202.150 50.495 -201.920 ;
        RECT 53.020 -202.020 60.830 -201.270 ;
        RECT 50.070 -202.470 50.390 -202.150 ;
        RECT 50.020 -202.750 50.460 -202.470 ;
        RECT 50.120 -203.360 50.390 -202.750 ;
        RECT 53.020 -203.320 53.220 -202.020 ;
        RECT 54.170 -202.040 60.830 -202.020 ;
        RECT 58.550 -202.060 60.830 -202.040 ;
        RECT 52.000 -203.360 53.220 -203.320 ;
        RECT 50.120 -203.740 53.220 -203.360 ;
        RECT 50.120 -204.260 50.390 -203.740 ;
        RECT 52.000 -203.790 53.220 -203.740 ;
        RECT 52.000 -203.800 53.200 -203.790 ;
        RECT 49.950 -204.610 50.470 -204.260 ;
        RECT 50.010 -204.900 50.410 -204.610 ;
        RECT 49.475 -205.130 50.475 -204.900 ;
        RECT 60.130 -215.750 60.830 -202.060 ;
        RECT 88.380 -202.550 88.700 -192.760 ;
        RECT 91.600 -202.550 92.540 -202.190 ;
        RECT 88.380 -202.840 92.540 -202.550 ;
        RECT 60.130 -215.800 62.950 -215.750 ;
        RECT 88.380 -215.800 88.700 -202.840 ;
        RECT 91.600 -203.150 92.540 -202.840 ;
        RECT 60.130 -216.640 88.740 -215.800 ;
        RECT 49.405 -217.450 50.405 -217.220 ;
        RECT 50.100 -217.700 50.350 -217.450 ;
        RECT 50.020 -218.070 50.430 -217.700 ;
        RECT 50.100 -218.360 50.350 -218.070 ;
        RECT 50.080 -218.810 53.160 -218.360 ;
        RECT 52.860 -221.560 53.060 -218.810 ;
        RECT 54.520 -221.500 55.210 -221.370 ;
        RECT 53.750 -221.550 56.120 -221.500 ;
        RECT 60.130 -221.550 60.830 -216.640 ;
        RECT 62.210 -216.810 88.740 -216.640 ;
        RECT 88.380 -216.960 88.700 -216.810 ;
        RECT 53.750 -221.560 60.830 -221.550 ;
        RECT 49.335 -222.440 50.335 -222.210 ;
        RECT 52.860 -222.310 60.830 -221.560 ;
        RECT 49.910 -222.760 50.230 -222.440 ;
        RECT 49.860 -223.040 50.300 -222.760 ;
        RECT 49.960 -223.650 50.230 -223.040 ;
        RECT 52.860 -223.610 53.060 -222.310 ;
        RECT 53.750 -222.340 60.830 -222.310 ;
        RECT 51.840 -223.650 53.060 -223.610 ;
        RECT 49.960 -224.030 53.060 -223.650 ;
        RECT 49.960 -224.550 50.230 -224.030 ;
        RECT 51.840 -224.080 53.060 -224.030 ;
        RECT 51.840 -224.090 53.040 -224.080 ;
        RECT 49.790 -224.900 50.310 -224.550 ;
        RECT 49.850 -225.190 50.250 -224.900 ;
        RECT 49.315 -225.420 50.315 -225.190 ;
        RECT 47.965 -237.220 48.965 -236.990 ;
        RECT 48.490 -237.460 48.910 -237.220 ;
        RECT 54.520 -237.460 55.210 -222.340 ;
        RECT 56.110 -222.440 60.830 -222.340 ;
        RECT 60.130 -222.460 60.830 -222.440 ;
        RECT 48.480 -237.540 55.210 -237.460 ;
        RECT 48.380 -237.840 55.210 -237.540 ;
        RECT 48.480 -237.860 55.210 -237.840 ;
        RECT 54.520 -237.970 55.210 -237.860 ;
      LAYER via ;
        RECT 89.610 176.460 89.950 176.810 ;
        RECT 83.150 166.260 83.490 166.670 ;
        RECT 51.100 156.410 51.460 156.950 ;
        RECT -233.120 -24.620 -232.580 -24.260 ;
        RECT -242.840 -56.650 -242.430 -56.310 ;
        RECT -253.060 -62.670 -252.800 -62.410 ;
        RECT 53.520 -182.840 53.880 -182.300 ;
        RECT 85.570 -192.560 85.910 -192.150 ;
        RECT 91.920 -202.820 92.180 -202.560 ;
      LAYER met2 ;
        RECT -390.150 -348.900 -380.150 326.100 ;
        RECT 89.570 177.180 90.520 326.090 ;
        RECT 89.330 176.370 90.520 177.180 ;
        RECT 89.330 176.200 90.290 176.370 ;
        RECT 50.830 166.880 84.170 166.930 ;
        RECT 50.740 165.690 84.170 166.880 ;
        RECT 50.740 157.860 51.560 165.690 ;
        RECT 51.000 157.230 51.520 157.860 ;
        RECT 50.770 155.930 51.910 157.230 ;
        RECT -243.050 -23.990 -234.030 -23.900 ;
        RECT -243.100 -24.160 -234.030 -23.990 ;
        RECT -233.400 -24.160 -232.100 -23.930 ;
        RECT -243.100 -24.680 -232.100 -24.160 ;
        RECT -243.100 -24.720 -234.030 -24.680 ;
        RECT -243.100 -57.330 -241.860 -24.720 ;
        RECT -233.400 -25.070 -232.100 -24.680 ;
        RECT -253.220 -62.820 -252.270 -62.350 ;
        RECT -252.750 -348.940 -252.270 -62.820 ;
        RECT 53.190 -183.120 54.330 -181.820 ;
        RECT 53.420 -183.750 53.940 -183.120 ;
        RECT 53.160 -191.580 53.980 -183.750 ;
        RECT 53.160 -192.770 86.590 -191.580 ;
        RECT 53.250 -192.820 86.590 -192.770 ;
        RECT 91.670 -202.240 92.480 -201.810 ;
        RECT 91.640 -203.090 92.500 -202.240 ;
        RECT 91.670 -203.510 92.480 -203.090 ;
        RECT 91.520 -348.870 92.480 -203.510 ;
        RECT 91.520 -348.900 92.330 -348.870 ;
        RECT 229.850 -348.900 239.850 326.100 ;
      LAYER via2 ;
        RECT -387.650 318.600 -382.650 323.600 ;
        RECT 89.760 316.660 90.210 325.600 ;
        RECT 232.350 318.600 237.350 323.600 ;
        RECT -387.650 -346.400 -382.650 -341.400 ;
        RECT -252.620 -348.540 -252.320 -339.530 ;
        RECT 91.740 -347.930 92.200 -339.980 ;
        RECT 232.350 -346.400 237.350 -341.400 ;
      LAYER met3 ;
        RECT -400.150 316.100 249.850 326.100 ;
        RECT -400.150 -348.900 249.850 -338.900 ;
    END
  END vccd1
  OBS
      LAYER li1 ;
        RECT 42.160 210.740 43.200 210.910 ;
        RECT 45.525 210.690 46.565 210.860 ;
        RECT 42.850 199.490 43.020 199.820 ;
        RECT 43.190 199.790 44.230 199.960 ;
        RECT 43.190 199.350 44.230 199.520 ;
        RECT 44.400 199.490 44.570 199.820 ;
        RECT 46.490 199.470 46.660 199.800 ;
        RECT 46.875 199.770 47.915 199.940 ;
        RECT 48.130 199.470 48.300 199.800 ;
        RECT 43.080 196.330 44.120 196.500 ;
        RECT 46.895 195.910 47.935 196.080 ;
        RECT 42.720 191.120 42.890 191.450 ;
        RECT 43.060 190.980 44.100 191.150 ;
        RECT 44.270 191.120 44.440 191.450 ;
        RECT 46.580 191.060 46.750 191.390 ;
        RECT 46.965 190.920 48.005 191.090 ;
        RECT 48.220 191.060 48.390 191.390 ;
        RECT 43.350 179.500 44.390 179.670 ;
        RECT 47.035 179.480 48.075 179.650 ;
        RECT 43.350 179.060 44.390 179.230 ;
        RECT 43.240 176.040 44.280 176.210 ;
        RECT 47.055 175.620 48.095 175.790 ;
        RECT 42.880 170.830 43.050 171.160 ;
        RECT 43.220 170.690 44.260 170.860 ;
        RECT 44.430 170.830 44.600 171.160 ;
        RECT 46.740 170.770 46.910 171.100 ;
        RECT 47.125 170.630 48.165 170.800 ;
        RECT 48.380 170.770 48.550 171.100 ;
        RECT -6.220 149.460 -6.050 149.790 ;
        RECT -5.880 149.320 -4.840 149.490 ;
        RECT -4.670 149.460 -4.500 149.790 ;
        RECT -1.920 149.420 -1.750 149.750 ;
        RECT -1.535 149.280 -0.495 149.450 ;
        RECT -0.280 149.420 -0.110 149.750 ;
        RECT 71.710 149.030 71.880 149.360 ;
        RECT 72.050 148.890 73.090 149.060 ;
        RECT 73.260 149.030 73.430 149.360 ;
        RECT 76.010 148.990 76.180 149.320 ;
        RECT 76.395 148.850 77.435 149.020 ;
        RECT 77.650 148.990 77.820 149.320 ;
        RECT -11.740 142.470 -11.570 142.970 ;
        RECT 8.810 142.470 8.980 142.970 ;
        RECT -11.400 142.240 8.640 142.410 ;
        RECT 66.190 142.040 66.360 142.540 ;
        RECT 86.740 142.040 86.910 142.540 ;
        RECT 66.530 141.810 86.570 141.980 ;
        RECT -11.400 137.160 8.640 137.330 ;
        RECT -11.740 136.600 -11.570 137.100 ;
        RECT 8.810 136.600 8.980 137.100 ;
        RECT 16.615 136.890 36.655 137.060 ;
        RECT 16.230 136.330 16.400 136.830 ;
        RECT 36.870 136.330 37.040 136.830 ;
        RECT 66.530 136.730 86.570 136.900 ;
        RECT 66.190 136.170 66.360 136.670 ;
        RECT 86.740 136.170 86.910 136.670 ;
        RECT 94.545 136.460 114.585 136.630 ;
        RECT 94.160 135.900 94.330 136.400 ;
        RECT 114.800 135.900 114.970 136.400 ;
        RECT -11.790 130.300 -11.620 130.800 ;
        RECT 8.760 130.300 8.930 130.800 ;
        RECT -11.450 130.070 8.590 130.240 ;
        RECT 16.290 130.140 16.460 130.640 ;
        RECT 36.930 130.140 37.100 130.640 ;
        RECT 16.675 129.910 36.715 130.080 ;
        RECT 66.140 129.870 66.310 130.370 ;
        RECT 86.690 129.870 86.860 130.370 ;
        RECT 66.480 129.640 86.520 129.810 ;
        RECT 94.220 129.710 94.390 130.210 ;
        RECT 114.860 129.710 115.030 130.210 ;
        RECT 94.605 129.480 114.645 129.650 ;
        RECT -11.660 125.040 8.380 125.210 ;
        RECT -12.000 124.480 -11.830 124.980 ;
        RECT 8.550 124.480 8.720 124.980 ;
        RECT 66.270 124.610 86.310 124.780 ;
        RECT 65.930 124.050 66.100 124.550 ;
        RECT 86.480 124.050 86.650 124.550 ;
        RECT 65.040 87.220 65.210 87.720 ;
        RECT 85.680 87.220 85.850 87.720 ;
        RECT 65.425 86.990 85.465 87.160 ;
        RECT -1.520 85.930 -1.350 86.430 ;
        RECT 19.120 85.930 19.290 86.430 ;
        RECT -1.135 85.700 18.905 85.870 ;
        RECT 65.230 84.130 85.270 84.300 ;
        RECT 64.890 83.570 65.060 84.070 ;
        RECT 85.440 83.570 85.610 84.070 ;
        RECT -1.330 82.840 18.710 83.010 ;
        RECT -1.670 82.280 -1.500 82.780 ;
        RECT 18.880 82.280 19.050 82.780 ;
        RECT 85.640 46.720 85.810 46.800 ;
        RECT 85.640 45.880 87.625 46.720 ;
        RECT 85.640 45.800 85.810 45.880 ;
        RECT 20.950 44.180 21.120 44.260 ;
        RECT 20.950 43.340 22.935 44.180 ;
        RECT 20.950 43.260 21.120 43.340 ;
        RECT 67.275 40.680 87.315 40.850 ;
        RECT 66.890 40.120 67.060 40.620 ;
        RECT 87.530 40.120 87.700 40.620 ;
        RECT 67.275 39.890 87.315 40.060 ;
        RECT -201.150 38.670 -200.650 38.840 ;
        RECT -219.140 38.410 -218.640 38.580 ;
        RECT -213.270 38.410 -212.770 38.580 ;
        RECT -206.970 38.460 -206.470 38.630 ;
        RECT -225.960 32.890 -225.630 33.060 ;
        RECT -225.660 31.680 -225.490 32.720 ;
        RECT -225.960 31.340 -225.630 31.510 ;
        RECT -225.920 28.590 -225.590 28.760 ;
        RECT -225.620 27.335 -225.450 28.375 ;
        RECT -225.920 26.950 -225.590 27.120 ;
        RECT -218.580 18.200 -218.410 38.240 ;
        RECT -213.500 18.200 -213.330 38.240 ;
        RECT -206.410 18.250 -206.240 38.290 ;
        RECT -201.380 18.460 -201.210 38.500 ;
        RECT 2.455 37.690 22.495 37.860 ;
        RECT 2.070 37.130 2.240 37.630 ;
        RECT 22.710 37.130 22.880 37.630 ;
        RECT 2.455 36.900 22.495 37.070 ;
        RECT 67.080 37.030 87.120 37.200 ;
        RECT 66.740 36.470 66.910 36.970 ;
        RECT 87.290 36.470 87.460 36.970 ;
        RECT 67.080 36.240 87.120 36.410 ;
        RECT 2.260 34.040 22.300 34.210 ;
        RECT 1.920 33.480 2.090 33.980 ;
        RECT 22.470 33.480 22.640 33.980 ;
        RECT 2.260 33.250 22.300 33.420 ;
        RECT -162.600 28.190 -162.100 28.360 ;
        RECT -158.950 28.340 -158.450 28.510 ;
        RECT -201.150 18.120 -200.650 18.290 ;
        RECT -219.140 17.860 -218.640 18.030 ;
        RECT -213.270 17.860 -212.770 18.030 ;
        RECT -206.970 17.910 -206.470 18.080 ;
        RECT -213.000 10.440 -212.500 10.610 ;
        RECT -206.810 10.380 -206.310 10.550 ;
        RECT -213.230 -9.815 -213.060 10.225 ;
        RECT -206.250 -9.875 -206.080 10.165 ;
        RECT -162.040 7.935 -161.870 27.975 ;
        RECT -159.180 8.130 -159.010 28.170 ;
        RECT -113.800 24.600 -113.300 24.770 ;
        RECT -110.150 24.750 -109.650 24.920 ;
        RECT -158.950 7.790 -158.450 7.960 ;
        RECT -162.600 7.550 -162.100 7.720 ;
        RECT -120.430 5.720 -119.430 5.890 ;
        RECT -120.350 3.905 -119.510 5.720 ;
        RECT -114.030 4.345 -113.860 24.385 ;
        RECT -113.240 4.345 -113.070 24.385 ;
        RECT -110.380 4.540 -110.210 24.580 ;
        RECT -109.590 4.540 -109.420 24.580 ;
        RECT 1.840 5.340 2.235 5.410 ;
        RECT -110.150 4.200 -109.650 4.370 ;
        RECT 1.840 4.340 2.240 5.340 ;
        RECT 3.440 4.340 3.840 5.440 ;
        RECT 5.920 5.360 6.315 5.430 ;
        RECT 5.920 4.360 6.320 5.360 ;
        RECT 7.520 4.360 7.920 5.460 ;
        RECT -113.800 3.960 -113.300 4.130 ;
        RECT 2.340 3.840 3.340 4.140 ;
        RECT 6.420 3.860 7.420 4.160 ;
        RECT 1.800 1.900 2.195 1.970 ;
        RECT 1.800 0.900 2.200 1.900 ;
        RECT 3.400 0.900 3.800 2.000 ;
        RECT 5.860 1.920 6.255 1.990 ;
        RECT 5.860 0.920 6.260 1.920 ;
        RECT 7.460 0.920 7.860 2.020 ;
        RECT 2.300 0.400 3.300 0.700 ;
        RECT 6.360 0.420 7.360 0.720 ;
        RECT -213.000 -10.200 -212.500 -10.030 ;
        RECT -206.810 -10.260 -206.310 -10.090 ;
        RECT -287.080 -16.360 -286.910 -15.320 ;
        RECT -275.990 -16.180 -275.660 -16.010 ;
        RECT -267.620 -16.050 -267.290 -15.880 ;
        RECT -247.330 -16.210 -247.000 -16.040 ;
        RECT -276.130 -17.390 -275.960 -16.350 ;
        RECT -275.690 -17.390 -275.520 -16.350 ;
        RECT -272.670 -17.280 -272.500 -16.240 ;
        RECT -267.320 -17.260 -267.150 -16.220 ;
        RECT -275.990 -17.730 -275.660 -17.560 ;
        RECT -267.620 -17.600 -267.290 -17.430 ;
        RECT -255.840 -17.550 -255.670 -16.510 ;
        RECT -255.400 -17.550 -255.230 -16.510 ;
        RECT -252.380 -17.440 -252.210 -16.400 ;
        RECT -247.030 -17.420 -246.860 -16.380 ;
        RECT -247.330 -17.760 -247.000 -17.590 ;
        RECT -287.030 -19.725 -286.860 -18.685 ;
        RECT -275.970 -19.820 -275.640 -19.650 ;
        RECT -267.560 -19.910 -267.230 -19.740 ;
        RECT -276.110 -21.075 -275.940 -20.035 ;
        RECT -272.250 -21.095 -272.080 -20.055 ;
        RECT -247.270 -20.070 -246.940 -19.900 ;
        RECT -267.260 -21.165 -267.090 -20.125 ;
        RECT -255.820 -21.235 -255.650 -20.195 ;
        RECT -251.960 -21.255 -251.790 -20.215 ;
        RECT -275.970 -21.460 -275.640 -21.290 ;
        RECT -246.970 -21.325 -246.800 -20.285 ;
        RECT -267.560 -21.550 -267.230 -21.380 ;
        RECT -247.270 -21.710 -246.940 -21.540 ;
        RECT -163.890 -38.370 -163.390 -38.200 ;
        RECT -160.240 -38.220 -159.740 -38.050 ;
        RECT -200.720 -39.260 -200.220 -39.090 ;
        RECT -218.710 -39.520 -218.210 -39.350 ;
        RECT -212.840 -39.520 -212.340 -39.350 ;
        RECT -206.540 -39.470 -206.040 -39.300 ;
        RECT -225.530 -45.040 -225.200 -44.870 ;
        RECT -225.230 -46.250 -225.060 -45.210 ;
        RECT -225.530 -46.590 -225.200 -46.420 ;
        RECT -225.490 -49.340 -225.160 -49.170 ;
        RECT -225.190 -50.595 -225.020 -49.555 ;
        RECT -225.490 -50.980 -225.160 -50.810 ;
        RECT -218.150 -59.730 -217.980 -39.690 ;
        RECT -213.070 -59.730 -212.900 -39.690 ;
        RECT -205.980 -59.680 -205.810 -39.640 ;
        RECT -200.950 -59.470 -200.780 -39.430 ;
        RECT -163.330 -58.625 -163.160 -38.585 ;
        RECT -160.470 -58.430 -160.300 -38.390 ;
        RECT -116.790 -40.220 -116.290 -40.050 ;
        RECT -113.140 -40.070 -112.640 -39.900 ;
        RECT -160.240 -58.770 -159.740 -58.600 ;
        RECT -163.890 -59.010 -163.390 -58.840 ;
        RECT -122.970 -58.970 -121.970 -58.800 ;
        RECT -200.720 -59.810 -200.220 -59.640 ;
        RECT -218.710 -60.070 -218.210 -59.900 ;
        RECT -212.840 -60.070 -212.340 -59.900 ;
        RECT -206.540 -60.020 -206.040 -59.850 ;
        RECT -122.890 -60.785 -122.050 -58.970 ;
        RECT -117.020 -60.475 -116.850 -40.435 ;
        RECT -116.230 -60.475 -116.060 -40.435 ;
        RECT -113.370 -60.280 -113.200 -40.240 ;
        RECT -112.580 -60.280 -112.410 -40.240 ;
        RECT 4.680 -59.310 24.720 -59.140 ;
        RECT 4.340 -59.870 4.510 -59.370 ;
        RECT 24.890 -59.870 25.060 -59.370 ;
        RECT 4.680 -60.100 24.720 -59.930 ;
        RECT -113.140 -60.620 -112.640 -60.450 ;
        RECT -116.790 -60.860 -116.290 -60.690 ;
        RECT 69.500 -62.300 89.540 -62.130 ;
        RECT 4.875 -62.960 24.915 -62.790 ;
        RECT 69.160 -62.860 69.330 -62.360 ;
        RECT 89.710 -62.860 89.880 -62.360 ;
        RECT 4.490 -63.520 4.660 -63.020 ;
        RECT 25.130 -63.520 25.300 -63.020 ;
        RECT 69.500 -63.090 89.540 -62.920 ;
        RECT 4.875 -63.750 24.915 -63.580 ;
        RECT 69.695 -65.950 89.735 -65.780 ;
        RECT 69.310 -66.510 69.480 -66.010 ;
        RECT 89.950 -66.510 90.120 -66.010 ;
        RECT 69.695 -66.740 89.735 -66.570 ;
        RECT -212.570 -67.490 -212.070 -67.320 ;
        RECT -206.380 -67.550 -205.880 -67.380 ;
        RECT -212.800 -87.745 -212.630 -67.705 ;
        RECT -205.820 -87.805 -205.650 -67.765 ;
        RECT 23.370 -69.230 23.540 -69.150 ;
        RECT 23.370 -70.070 25.355 -69.230 ;
        RECT 23.370 -70.150 23.540 -70.070 ;
        RECT 88.060 -71.770 88.230 -71.690 ;
        RECT 88.060 -72.610 90.045 -71.770 ;
        RECT 88.060 -72.690 88.230 -72.610 ;
        RECT -212.570 -88.130 -212.070 -87.960 ;
        RECT -206.380 -88.190 -205.880 -88.020 ;
        RECT 0.750 -108.670 0.920 -108.170 ;
        RECT 21.300 -108.670 21.470 -108.170 ;
        RECT 1.090 -108.900 21.130 -108.730 ;
        RECT 67.310 -109.960 67.480 -109.460 ;
        RECT 87.860 -109.960 88.030 -109.460 ;
        RECT 67.650 -110.190 87.690 -110.020 ;
        RECT 1.285 -111.760 21.325 -111.590 ;
        RECT 0.900 -112.320 1.070 -111.820 ;
        RECT 21.540 -112.320 21.710 -111.820 ;
        RECT 67.845 -113.050 87.885 -112.880 ;
        RECT 67.460 -113.610 67.630 -113.110 ;
        RECT 88.100 -113.610 88.270 -113.110 ;
        RECT -9.580 -150.870 -9.410 -150.370 ;
        RECT 10.970 -150.870 11.140 -150.370 ;
        RECT 68.350 -150.440 68.520 -149.940 ;
        RECT 88.900 -150.440 89.070 -149.940 ;
        RECT 68.690 -150.670 88.730 -150.500 ;
        RECT -9.240 -151.100 10.800 -150.930 ;
        RECT 68.900 -155.700 88.940 -155.530 ;
        RECT 97.025 -155.540 117.065 -155.370 ;
        RECT -9.030 -156.130 11.010 -155.960 ;
        RECT 19.095 -155.970 39.135 -155.800 ;
        RECT -9.370 -156.690 -9.200 -156.190 ;
        RECT 11.180 -156.690 11.350 -156.190 ;
        RECT 18.710 -156.530 18.880 -156.030 ;
        RECT 39.350 -156.530 39.520 -156.030 ;
        RECT 68.560 -156.260 68.730 -155.760 ;
        RECT 89.110 -156.260 89.280 -155.760 ;
        RECT 96.640 -156.100 96.810 -155.600 ;
        RECT 117.280 -156.100 117.450 -155.600 ;
        RECT -9.320 -162.990 -9.150 -162.490 ;
        RECT 11.230 -162.990 11.400 -162.490 ;
        RECT 18.650 -162.720 18.820 -162.220 ;
        RECT 39.290 -162.720 39.460 -162.220 ;
        RECT 68.610 -162.560 68.780 -162.060 ;
        RECT 89.160 -162.560 89.330 -162.060 ;
        RECT 96.580 -162.290 96.750 -161.790 ;
        RECT 117.220 -162.290 117.390 -161.790 ;
        RECT 96.965 -162.520 117.005 -162.350 ;
        RECT 19.035 -162.950 39.075 -162.780 ;
        RECT 68.950 -162.790 88.990 -162.620 ;
        RECT -8.980 -163.220 11.060 -163.050 ;
        RECT 68.950 -167.870 88.990 -167.700 ;
        RECT -8.980 -168.300 11.060 -168.130 ;
        RECT -9.320 -168.860 -9.150 -168.360 ;
        RECT 11.230 -168.860 11.400 -168.360 ;
        RECT 68.610 -168.430 68.780 -167.930 ;
        RECT 89.160 -168.430 89.330 -167.930 ;
        RECT -3.800 -175.680 -3.630 -175.350 ;
        RECT -3.460 -175.380 -2.420 -175.210 ;
        RECT -2.250 -175.680 -2.080 -175.350 ;
        RECT 0.500 -175.640 0.670 -175.310 ;
        RECT 0.885 -175.340 1.925 -175.170 ;
        RECT 74.130 -175.250 74.300 -174.920 ;
        RECT 74.470 -174.950 75.510 -174.780 ;
        RECT 75.680 -175.250 75.850 -174.920 ;
        RECT 78.430 -175.210 78.600 -174.880 ;
        RECT 78.815 -174.910 79.855 -174.740 ;
        RECT 80.070 -175.210 80.240 -174.880 ;
        RECT 2.140 -175.640 2.310 -175.310 ;
        RECT 45.300 -197.050 45.470 -196.720 ;
        RECT 45.640 -196.750 46.680 -196.580 ;
        RECT 46.850 -197.050 47.020 -196.720 ;
        RECT 49.160 -196.990 49.330 -196.660 ;
        RECT 49.545 -196.690 50.585 -196.520 ;
        RECT 50.800 -196.990 50.970 -196.660 ;
        RECT 49.475 -201.680 50.515 -201.510 ;
        RECT 45.660 -202.100 46.700 -201.930 ;
        RECT 45.770 -205.120 46.810 -204.950 ;
        RECT 45.770 -205.560 46.810 -205.390 ;
        RECT 49.455 -205.540 50.495 -205.370 ;
        RECT 45.140 -217.340 45.310 -217.010 ;
        RECT 45.480 -217.040 46.520 -216.870 ;
        RECT 46.690 -217.340 46.860 -217.010 ;
        RECT 49.000 -217.280 49.170 -216.950 ;
        RECT 49.385 -216.980 50.425 -216.810 ;
        RECT 50.640 -217.280 50.810 -216.950 ;
        RECT 49.315 -221.970 50.355 -221.800 ;
        RECT 45.500 -222.390 46.540 -222.220 ;
        RECT 45.270 -225.710 45.440 -225.380 ;
        RECT 45.610 -225.410 46.650 -225.240 ;
        RECT 45.610 -225.850 46.650 -225.680 ;
        RECT 46.820 -225.710 46.990 -225.380 ;
        RECT 48.910 -225.690 49.080 -225.360 ;
        RECT 49.295 -225.830 50.335 -225.660 ;
        RECT 50.550 -225.690 50.720 -225.360 ;
        RECT 44.580 -236.800 45.620 -236.630 ;
        RECT 47.945 -236.750 48.985 -236.580 ;
      LAYER mcon ;
        RECT 42.240 210.740 43.120 210.910 ;
        RECT 45.605 210.690 46.485 210.860 ;
        RECT 43.270 199.790 44.150 199.960 ;
        RECT 42.850 199.570 43.020 199.740 ;
        RECT 44.400 199.570 44.570 199.740 ;
        RECT 43.270 199.350 44.150 199.520 ;
        RECT 46.955 199.770 47.835 199.940 ;
        RECT 46.490 199.550 46.660 199.720 ;
        RECT 48.130 199.550 48.300 199.720 ;
        RECT 43.160 196.330 44.040 196.500 ;
        RECT 46.975 195.910 47.855 196.080 ;
        RECT 42.720 191.200 42.890 191.370 ;
        RECT 44.270 191.200 44.440 191.370 ;
        RECT 43.140 190.980 44.020 191.150 ;
        RECT 46.580 191.140 46.750 191.310 ;
        RECT 48.220 191.140 48.390 191.310 ;
        RECT 47.045 190.920 47.925 191.090 ;
        RECT 43.430 179.500 44.310 179.670 ;
        RECT 47.115 179.480 47.995 179.650 ;
        RECT 43.430 179.060 44.310 179.230 ;
        RECT 43.320 176.040 44.200 176.210 ;
        RECT 47.135 175.620 48.015 175.790 ;
        RECT 42.880 170.910 43.050 171.080 ;
        RECT 44.430 170.910 44.600 171.080 ;
        RECT 43.300 170.690 44.180 170.860 ;
        RECT 46.740 170.850 46.910 171.020 ;
        RECT 48.380 170.850 48.550 171.020 ;
        RECT 47.205 170.630 48.085 170.800 ;
        RECT -6.220 149.540 -6.050 149.710 ;
        RECT -4.670 149.540 -4.500 149.710 ;
        RECT -5.800 149.320 -4.920 149.490 ;
        RECT -1.920 149.500 -1.750 149.670 ;
        RECT -0.280 149.500 -0.110 149.670 ;
        RECT -1.455 149.280 -0.575 149.450 ;
        RECT 71.710 149.110 71.880 149.280 ;
        RECT 73.260 149.110 73.430 149.280 ;
        RECT 72.130 148.890 73.010 149.060 ;
        RECT 76.010 149.070 76.180 149.240 ;
        RECT 77.650 149.070 77.820 149.240 ;
        RECT 76.475 148.850 77.355 149.020 ;
        RECT -11.740 142.550 -11.570 142.890 ;
        RECT 8.810 142.550 8.980 142.890 ;
        RECT -11.320 142.240 8.560 142.410 ;
        RECT 66.190 142.120 66.360 142.460 ;
        RECT 86.740 142.120 86.910 142.460 ;
        RECT 66.610 141.810 86.490 141.980 ;
        RECT -11.320 137.160 8.560 137.330 ;
        RECT -11.740 136.680 -11.570 137.020 ;
        RECT 8.810 136.680 8.980 137.020 ;
        RECT 16.695 136.890 36.575 137.060 ;
        RECT 16.230 136.410 16.400 136.750 ;
        RECT 36.870 136.410 37.040 136.750 ;
        RECT 66.610 136.730 86.490 136.900 ;
        RECT 66.190 136.250 66.360 136.590 ;
        RECT 86.740 136.250 86.910 136.590 ;
        RECT 94.625 136.460 114.505 136.630 ;
        RECT 94.160 135.980 94.330 136.320 ;
        RECT 114.800 135.980 114.970 136.320 ;
        RECT -11.790 130.380 -11.620 130.720 ;
        RECT 8.760 130.380 8.930 130.720 ;
        RECT -11.370 130.070 8.510 130.240 ;
        RECT 16.290 130.220 16.460 130.560 ;
        RECT 36.930 130.220 37.100 130.560 ;
        RECT 16.755 129.910 36.635 130.080 ;
        RECT 66.140 129.950 66.310 130.290 ;
        RECT 86.690 129.950 86.860 130.290 ;
        RECT 66.560 129.640 86.440 129.810 ;
        RECT 94.220 129.790 94.390 130.130 ;
        RECT 114.860 129.790 115.030 130.130 ;
        RECT 94.685 129.480 114.565 129.650 ;
        RECT -11.580 125.040 8.300 125.210 ;
        RECT -12.000 124.560 -11.830 124.900 ;
        RECT 8.550 124.560 8.720 124.900 ;
        RECT 66.350 124.610 86.230 124.780 ;
        RECT 65.930 124.130 66.100 124.470 ;
        RECT 86.480 124.130 86.650 124.470 ;
        RECT 65.040 87.300 65.210 87.640 ;
        RECT 85.680 87.300 85.850 87.640 ;
        RECT 65.505 86.990 85.385 87.160 ;
        RECT -1.520 86.010 -1.350 86.350 ;
        RECT 19.120 86.010 19.290 86.350 ;
        RECT -1.055 85.700 18.825 85.870 ;
        RECT 65.310 84.130 85.190 84.300 ;
        RECT 64.890 83.650 65.060 83.990 ;
        RECT 85.440 83.650 85.610 83.990 ;
        RECT -1.250 82.840 18.630 83.010 ;
        RECT -1.670 82.360 -1.500 82.700 ;
        RECT 18.880 82.360 19.050 82.700 ;
        RECT 85.640 45.880 87.625 46.720 ;
        RECT 20.950 43.340 22.935 44.180 ;
        RECT 67.355 40.680 87.235 40.850 ;
        RECT 66.890 40.200 67.060 40.540 ;
        RECT 87.530 40.200 87.700 40.540 ;
        RECT 67.355 39.890 87.235 40.060 ;
        RECT -201.070 38.670 -200.730 38.840 ;
        RECT -219.060 38.410 -218.720 38.580 ;
        RECT -213.190 38.410 -212.850 38.580 ;
        RECT -206.890 38.460 -206.550 38.630 ;
        RECT -225.880 32.890 -225.710 33.060 ;
        RECT -225.660 31.760 -225.490 32.640 ;
        RECT -225.880 31.340 -225.710 31.510 ;
        RECT -225.840 28.590 -225.670 28.760 ;
        RECT -225.620 27.415 -225.450 28.295 ;
        RECT -225.840 26.950 -225.670 27.120 ;
        RECT -218.580 18.280 -218.410 38.160 ;
        RECT -213.500 18.280 -213.330 38.160 ;
        RECT -206.410 18.330 -206.240 38.210 ;
        RECT -201.380 18.540 -201.210 38.420 ;
        RECT 2.535 37.690 22.415 37.860 ;
        RECT 2.070 37.210 2.240 37.550 ;
        RECT 22.710 37.210 22.880 37.550 ;
        RECT 2.535 36.900 22.415 37.070 ;
        RECT 67.160 37.030 87.040 37.200 ;
        RECT 66.740 36.550 66.910 36.890 ;
        RECT 87.290 36.550 87.460 36.890 ;
        RECT 67.160 36.240 87.040 36.410 ;
        RECT 2.340 34.040 22.220 34.210 ;
        RECT 1.920 33.560 2.090 33.900 ;
        RECT 22.470 33.560 22.640 33.900 ;
        RECT 2.340 33.250 22.220 33.420 ;
        RECT -162.520 28.190 -162.180 28.360 ;
        RECT -158.870 28.340 -158.530 28.510 ;
        RECT -201.070 18.120 -200.730 18.290 ;
        RECT -219.060 17.860 -218.720 18.030 ;
        RECT -213.190 17.860 -212.850 18.030 ;
        RECT -206.890 17.910 -206.550 18.080 ;
        RECT -212.920 10.440 -212.580 10.610 ;
        RECT -206.730 10.380 -206.390 10.550 ;
        RECT -213.230 -9.735 -213.060 10.145 ;
        RECT -206.250 -9.795 -206.080 10.085 ;
        RECT -162.040 8.015 -161.870 27.895 ;
        RECT -159.180 8.210 -159.010 28.090 ;
        RECT -113.720 24.600 -113.380 24.770 ;
        RECT -110.070 24.750 -109.730 24.920 ;
        RECT -158.870 7.790 -158.530 7.960 ;
        RECT -162.520 7.550 -162.180 7.720 ;
        RECT -114.030 4.425 -113.860 24.305 ;
        RECT -113.240 4.425 -113.070 24.305 ;
        RECT -110.380 4.620 -110.210 24.500 ;
        RECT -109.590 4.620 -109.420 24.500 ;
        RECT 1.940 4.540 2.140 5.240 ;
        RECT -110.070 4.200 -109.730 4.370 ;
        RECT 3.540 4.540 3.740 5.240 ;
        RECT 6.020 4.560 6.220 5.260 ;
        RECT 7.620 4.560 7.820 5.260 ;
        RECT -113.720 3.960 -113.380 4.130 ;
        RECT 2.440 3.940 3.240 4.110 ;
        RECT 6.520 3.960 7.320 4.130 ;
        RECT 1.900 1.100 2.100 1.800 ;
        RECT 3.500 1.100 3.700 1.800 ;
        RECT 5.960 1.120 6.160 1.820 ;
        RECT 7.560 1.120 7.760 1.820 ;
        RECT 2.400 0.500 3.200 0.670 ;
        RECT 6.460 0.520 7.260 0.690 ;
        RECT -212.920 -10.200 -212.580 -10.030 ;
        RECT -206.730 -10.260 -206.390 -10.090 ;
        RECT -287.080 -16.280 -286.910 -15.400 ;
        RECT -275.910 -16.180 -275.740 -16.010 ;
        RECT -267.540 -16.050 -267.370 -15.880 ;
        RECT -247.250 -16.210 -247.080 -16.040 ;
        RECT -276.130 -17.310 -275.960 -16.430 ;
        RECT -275.690 -17.310 -275.520 -16.430 ;
        RECT -272.670 -17.200 -272.500 -16.320 ;
        RECT -267.320 -17.180 -267.150 -16.300 ;
        RECT -275.910 -17.730 -275.740 -17.560 ;
        RECT -267.540 -17.600 -267.370 -17.430 ;
        RECT -255.840 -17.470 -255.670 -16.590 ;
        RECT -255.400 -17.470 -255.230 -16.590 ;
        RECT -252.380 -17.360 -252.210 -16.480 ;
        RECT -247.030 -17.340 -246.860 -16.460 ;
        RECT -247.250 -17.760 -247.080 -17.590 ;
        RECT -287.030 -19.645 -286.860 -18.765 ;
        RECT -275.890 -19.820 -275.720 -19.650 ;
        RECT -267.480 -19.910 -267.310 -19.740 ;
        RECT -276.110 -20.995 -275.940 -20.115 ;
        RECT -247.190 -20.070 -247.020 -19.900 ;
        RECT -272.250 -21.015 -272.080 -20.135 ;
        RECT -267.260 -21.085 -267.090 -20.205 ;
        RECT -255.820 -21.155 -255.650 -20.275 ;
        RECT -251.960 -21.175 -251.790 -20.295 ;
        RECT -246.970 -21.245 -246.800 -20.365 ;
        RECT -275.890 -21.460 -275.720 -21.290 ;
        RECT -267.480 -21.550 -267.310 -21.380 ;
        RECT -247.190 -21.710 -247.020 -21.540 ;
        RECT -163.810 -38.370 -163.470 -38.200 ;
        RECT -160.160 -38.220 -159.820 -38.050 ;
        RECT -200.640 -39.260 -200.300 -39.090 ;
        RECT -218.630 -39.520 -218.290 -39.350 ;
        RECT -212.760 -39.520 -212.420 -39.350 ;
        RECT -206.460 -39.470 -206.120 -39.300 ;
        RECT -225.450 -45.040 -225.280 -44.870 ;
        RECT -225.230 -46.170 -225.060 -45.290 ;
        RECT -225.450 -46.590 -225.280 -46.420 ;
        RECT -225.410 -49.340 -225.240 -49.170 ;
        RECT -225.190 -50.515 -225.020 -49.635 ;
        RECT -225.410 -50.980 -225.240 -50.810 ;
        RECT -218.150 -59.650 -217.980 -39.770 ;
        RECT -213.070 -59.650 -212.900 -39.770 ;
        RECT -205.980 -59.600 -205.810 -39.720 ;
        RECT -200.950 -59.390 -200.780 -39.510 ;
        RECT -163.330 -58.545 -163.160 -38.665 ;
        RECT -160.470 -58.350 -160.300 -38.470 ;
        RECT -116.710 -40.220 -116.370 -40.050 ;
        RECT -113.060 -40.070 -112.720 -39.900 ;
        RECT -160.160 -58.770 -159.820 -58.600 ;
        RECT -163.810 -59.010 -163.470 -58.840 ;
        RECT -200.640 -59.810 -200.300 -59.640 ;
        RECT -218.630 -60.070 -218.290 -59.900 ;
        RECT -212.760 -60.070 -212.420 -59.900 ;
        RECT -206.460 -60.020 -206.120 -59.850 ;
        RECT -117.020 -60.395 -116.850 -40.515 ;
        RECT -116.230 -60.395 -116.060 -40.515 ;
        RECT -113.370 -60.200 -113.200 -40.320 ;
        RECT -112.580 -60.200 -112.410 -40.320 ;
        RECT 4.760 -59.310 24.640 -59.140 ;
        RECT 4.340 -59.790 4.510 -59.450 ;
        RECT 24.890 -59.790 25.060 -59.450 ;
        RECT 4.760 -60.100 24.640 -59.930 ;
        RECT -113.060 -60.620 -112.720 -60.450 ;
        RECT -116.710 -60.860 -116.370 -60.690 ;
        RECT 69.580 -62.300 89.460 -62.130 ;
        RECT 69.160 -62.780 69.330 -62.440 ;
        RECT 4.955 -62.960 24.835 -62.790 ;
        RECT 89.710 -62.780 89.880 -62.440 ;
        RECT 4.490 -63.440 4.660 -63.100 ;
        RECT 69.580 -63.090 89.460 -62.920 ;
        RECT 25.130 -63.440 25.300 -63.100 ;
        RECT 4.955 -63.750 24.835 -63.580 ;
        RECT 69.775 -65.950 89.655 -65.780 ;
        RECT 69.310 -66.430 69.480 -66.090 ;
        RECT 89.950 -66.430 90.120 -66.090 ;
        RECT 69.775 -66.740 89.655 -66.570 ;
        RECT -212.490 -67.490 -212.150 -67.320 ;
        RECT -206.300 -67.550 -205.960 -67.380 ;
        RECT -212.800 -87.665 -212.630 -67.785 ;
        RECT -205.820 -87.725 -205.650 -67.845 ;
        RECT 23.370 -70.070 25.355 -69.230 ;
        RECT 88.060 -72.610 90.045 -71.770 ;
        RECT -212.490 -88.130 -212.150 -87.960 ;
        RECT -206.300 -88.190 -205.960 -88.020 ;
        RECT 0.750 -108.590 0.920 -108.250 ;
        RECT 21.300 -108.590 21.470 -108.250 ;
        RECT 1.170 -108.900 21.050 -108.730 ;
        RECT 67.310 -109.880 67.480 -109.540 ;
        RECT 87.860 -109.880 88.030 -109.540 ;
        RECT 67.730 -110.190 87.610 -110.020 ;
        RECT 1.365 -111.760 21.245 -111.590 ;
        RECT 0.900 -112.240 1.070 -111.900 ;
        RECT 21.540 -112.240 21.710 -111.900 ;
        RECT 67.925 -113.050 87.805 -112.880 ;
        RECT 67.460 -113.530 67.630 -113.190 ;
        RECT 88.100 -113.530 88.270 -113.190 ;
        RECT 68.350 -150.360 68.520 -150.020 ;
        RECT -9.580 -150.790 -9.410 -150.450 ;
        RECT 88.900 -150.360 89.070 -150.020 ;
        RECT 10.970 -150.790 11.140 -150.450 ;
        RECT 68.770 -150.670 88.650 -150.500 ;
        RECT -9.160 -151.100 10.720 -150.930 ;
        RECT 68.980 -155.700 88.860 -155.530 ;
        RECT 97.105 -155.540 116.985 -155.370 ;
        RECT -8.950 -156.130 10.930 -155.960 ;
        RECT 19.175 -155.970 39.055 -155.800 ;
        RECT -9.370 -156.610 -9.200 -156.270 ;
        RECT 11.180 -156.610 11.350 -156.270 ;
        RECT 18.710 -156.450 18.880 -156.110 ;
        RECT 39.350 -156.450 39.520 -156.110 ;
        RECT 68.560 -156.180 68.730 -155.840 ;
        RECT 89.110 -156.180 89.280 -155.840 ;
        RECT 96.640 -156.020 96.810 -155.680 ;
        RECT 117.280 -156.020 117.450 -155.680 ;
        RECT -9.320 -162.910 -9.150 -162.570 ;
        RECT 11.230 -162.910 11.400 -162.570 ;
        RECT 18.650 -162.640 18.820 -162.300 ;
        RECT 39.290 -162.640 39.460 -162.300 ;
        RECT 68.610 -162.480 68.780 -162.140 ;
        RECT 89.160 -162.480 89.330 -162.140 ;
        RECT 96.580 -162.210 96.750 -161.870 ;
        RECT 117.220 -162.210 117.390 -161.870 ;
        RECT 97.045 -162.520 116.925 -162.350 ;
        RECT 19.115 -162.950 38.995 -162.780 ;
        RECT 69.030 -162.790 88.910 -162.620 ;
        RECT -8.900 -163.220 10.980 -163.050 ;
        RECT 69.030 -167.870 88.910 -167.700 ;
        RECT -8.900 -168.300 10.980 -168.130 ;
        RECT 68.610 -168.350 68.780 -168.010 ;
        RECT -9.320 -168.780 -9.150 -168.440 ;
        RECT 89.160 -168.350 89.330 -168.010 ;
        RECT 11.230 -168.780 11.400 -168.440 ;
        RECT 74.550 -174.950 75.430 -174.780 ;
        RECT 74.130 -175.170 74.300 -175.000 ;
        RECT -3.380 -175.380 -2.500 -175.210 ;
        RECT -3.800 -175.600 -3.630 -175.430 ;
        RECT -2.250 -175.600 -2.080 -175.430 ;
        RECT 0.965 -175.340 1.845 -175.170 ;
        RECT 75.680 -175.170 75.850 -175.000 ;
        RECT 78.895 -174.910 79.775 -174.740 ;
        RECT 78.430 -175.130 78.600 -174.960 ;
        RECT 80.070 -175.130 80.240 -174.960 ;
        RECT 0.500 -175.560 0.670 -175.390 ;
        RECT 2.140 -175.560 2.310 -175.390 ;
        RECT 45.720 -196.750 46.600 -196.580 ;
        RECT 45.300 -196.970 45.470 -196.800 ;
        RECT 46.850 -196.970 47.020 -196.800 ;
        RECT 49.625 -196.690 50.505 -196.520 ;
        RECT 49.160 -196.910 49.330 -196.740 ;
        RECT 50.800 -196.910 50.970 -196.740 ;
        RECT 49.555 -201.680 50.435 -201.510 ;
        RECT 45.740 -202.100 46.620 -201.930 ;
        RECT 45.850 -205.120 46.730 -204.950 ;
        RECT 45.850 -205.560 46.730 -205.390 ;
        RECT 49.535 -205.540 50.415 -205.370 ;
        RECT 45.560 -217.040 46.440 -216.870 ;
        RECT 45.140 -217.260 45.310 -217.090 ;
        RECT 46.690 -217.260 46.860 -217.090 ;
        RECT 49.465 -216.980 50.345 -216.810 ;
        RECT 49.000 -217.200 49.170 -217.030 ;
        RECT 50.640 -217.200 50.810 -217.030 ;
        RECT 49.395 -221.970 50.275 -221.800 ;
        RECT 45.580 -222.390 46.460 -222.220 ;
        RECT 45.690 -225.410 46.570 -225.240 ;
        RECT 45.270 -225.630 45.440 -225.460 ;
        RECT 46.820 -225.630 46.990 -225.460 ;
        RECT 45.690 -225.850 46.570 -225.680 ;
        RECT 48.910 -225.610 49.080 -225.440 ;
        RECT 50.550 -225.610 50.720 -225.440 ;
        RECT 49.375 -225.830 50.255 -225.660 ;
        RECT 44.660 -236.800 45.540 -236.630 ;
        RECT 48.025 -236.750 48.905 -236.580 ;
      LAYER met1 ;
        RECT 42.180 210.710 43.180 210.940 ;
        RECT 42.810 209.320 43.080 210.710 ;
        RECT 45.545 210.660 46.545 210.890 ;
        RECT 45.820 209.320 46.080 210.660 ;
        RECT 42.810 209.090 46.080 209.320 ;
        RECT 44.500 204.980 44.780 209.090 ;
        RECT 44.500 204.540 45.740 204.980 ;
        RECT 45.170 203.740 45.720 204.540 ;
        RECT 42.780 203.190 48.430 203.740 ;
        RECT 42.780 202.530 43.030 203.190 ;
        RECT 42.780 202.030 43.040 202.530 ;
        RECT 42.790 199.820 43.040 202.030 ;
        RECT 45.320 202.020 45.590 202.060 ;
        RECT 45.320 201.990 47.160 202.020 ;
        RECT 45.320 201.750 47.180 201.990 ;
        RECT 43.820 201.260 44.080 201.270 ;
        RECT 45.320 201.260 45.590 201.750 ;
        RECT 43.820 200.900 45.590 201.260 ;
        RECT 43.820 199.990 44.080 200.900 ;
        RECT 45.320 200.060 45.590 200.900 ;
        RECT 42.750 199.800 43.040 199.820 ;
        RECT 42.750 199.510 43.050 199.800 ;
        RECT 43.210 199.760 44.210 199.990 ;
        RECT 42.750 199.490 43.040 199.510 ;
        RECT 43.210 199.320 44.210 199.550 ;
        RECT 44.360 199.490 44.640 199.820 ;
        RECT 43.650 196.530 43.940 199.320 ;
        RECT 45.320 198.380 45.630 200.060 ;
        RECT 47.040 199.970 47.180 201.750 ;
        RECT 46.400 199.780 46.680 199.790 ;
        RECT 46.400 199.490 46.690 199.780 ;
        RECT 46.895 199.740 47.895 199.970 ;
        RECT 48.110 199.790 48.420 203.190 ;
        RECT 46.400 199.460 46.680 199.490 ;
        RECT 48.080 199.460 48.420 199.790 ;
        RECT 48.110 199.450 48.420 199.460 ;
        RECT 45.320 197.440 46.140 198.380 ;
        RECT 45.320 196.690 45.630 197.440 ;
        RECT 43.100 196.300 44.100 196.530 ;
        RECT 45.360 195.000 45.630 196.690 ;
        RECT 46.915 195.880 47.915 196.110 ;
        RECT 47.100 195.000 47.320 195.880 ;
        RECT 45.360 194.700 47.320 195.000 ;
        RECT 45.360 194.690 45.630 194.700 ;
        RECT 42.640 191.120 42.920 191.450 ;
        RECT 43.080 190.950 44.080 191.180 ;
        RECT 44.230 190.980 44.610 191.540 ;
        RECT 46.450 190.990 46.790 191.490 ;
        RECT 43.630 189.450 43.960 190.950 ;
        RECT 46.985 190.890 47.985 191.120 ;
        RECT 48.180 191.060 48.460 191.390 ;
        RECT 47.010 189.450 47.340 190.890 ;
        RECT 43.630 189.300 47.340 189.450 ;
        RECT 43.670 189.220 47.340 189.300 ;
        RECT 45.250 187.810 46.490 189.220 ;
        RECT 45.480 181.730 45.750 181.770 ;
        RECT 45.480 181.700 47.320 181.730 ;
        RECT 45.480 181.460 47.340 181.700 ;
        RECT 43.980 180.970 44.240 180.980 ;
        RECT 45.480 180.970 45.750 181.460 ;
        RECT 43.980 180.610 45.750 180.970 ;
        RECT 43.980 179.700 44.240 180.610 ;
        RECT 45.480 179.770 45.750 180.610 ;
        RECT 43.370 179.470 44.370 179.700 ;
        RECT 43.370 179.030 44.370 179.260 ;
        RECT 43.810 176.240 44.100 179.030 ;
        RECT 45.480 178.090 45.790 179.770 ;
        RECT 47.200 179.680 47.340 181.460 ;
        RECT 47.055 179.450 48.055 179.680 ;
        RECT 45.480 177.150 46.300 178.090 ;
        RECT 45.480 176.400 45.790 177.150 ;
        RECT 43.260 176.010 44.260 176.240 ;
        RECT 45.520 174.710 45.790 176.400 ;
        RECT 47.075 175.590 48.075 175.820 ;
        RECT 47.260 174.710 47.480 175.590 ;
        RECT 45.520 174.410 47.480 174.710 ;
        RECT 45.520 174.400 45.790 174.410 ;
        RECT 42.800 170.830 43.080 171.160 ;
        RECT 43.240 170.660 44.240 170.890 ;
        RECT 44.390 170.690 44.770 171.250 ;
        RECT 46.610 170.700 46.950 171.200 ;
        RECT 43.790 169.160 44.120 170.660 ;
        RECT 47.145 170.600 48.145 170.830 ;
        RECT 48.340 170.770 48.620 171.100 ;
        RECT 47.170 169.160 47.500 170.600 ;
        RECT 43.790 169.010 47.500 169.160 ;
        RECT 43.830 168.930 47.500 169.010 ;
        RECT 31.010 162.120 34.080 166.160 ;
        RECT 44.880 163.420 46.290 168.930 ;
        RECT 44.880 163.280 75.010 163.420 ;
        RECT 44.880 162.590 75.020 163.280 ;
        RECT 44.880 162.530 46.290 162.590 ;
        RECT 31.270 160.790 33.540 162.120 ;
        RECT 31.270 160.150 33.710 160.790 ;
        RECT 33.080 157.690 33.710 160.150 ;
        RECT -3.330 156.850 33.740 157.690 ;
        RECT -17.710 151.800 -14.750 151.810 ;
        RECT -3.290 151.800 -2.960 156.850 ;
        RECT -17.710 151.770 -2.960 151.800 ;
        RECT -17.710 151.500 -2.970 151.770 ;
        RECT 74.730 151.550 75.020 162.590 ;
        RECT -17.710 151.490 -14.750 151.500 ;
        RECT -17.660 124.990 -17.050 151.490 ;
        RECT -3.220 151.240 -2.970 151.500 ;
        RECT 74.710 151.430 75.020 151.550 ;
        RECT -4.740 151.220 -4.600 151.230 ;
        RECT -3.470 151.220 -2.970 151.240 ;
        RECT 60.220 151.370 63.180 151.380 ;
        RECT 74.710 151.370 74.960 151.430 ;
        RECT -4.740 151.190 -1.700 151.220 ;
        RECT -4.740 150.990 -1.690 151.190 ;
        RECT 60.220 151.070 74.960 151.370 ;
        RECT 60.220 151.060 63.180 151.070 ;
        RECT -4.720 150.800 -1.690 150.990 ;
        RECT -6.250 149.430 -6.010 149.820 ;
        RECT -4.720 149.770 -4.480 150.800 ;
        RECT -5.860 149.290 -4.860 149.520 ;
        RECT -4.720 149.480 -4.470 149.770 ;
        RECT -4.720 149.390 -4.480 149.480 ;
        RECT -5.850 149.190 -4.860 149.290 ;
        RECT -16.690 146.250 -16.010 146.290 ;
        RECT -14.060 146.250 -13.590 146.310 ;
        RECT -16.690 145.660 -13.590 146.250 ;
        RECT -3.470 146.180 -3.190 150.800 ;
        RECT -1.950 149.370 -1.690 150.800 ;
        RECT -0.280 149.730 -0.080 149.770 ;
        RECT -1.510 149.480 -0.470 149.490 ;
        RECT -1.515 149.250 -0.470 149.480 ;
        RECT -0.310 149.440 -0.080 149.730 ;
        RECT -0.280 149.380 -0.080 149.440 ;
        RECT -1.510 149.160 -0.470 149.250 ;
        RECT -1.470 149.150 -0.470 149.160 ;
        RECT -11.620 145.700 -3.190 146.180 ;
        RECT -11.620 145.690 -3.460 145.700 ;
        RECT -11.530 145.680 -3.490 145.690 ;
        RECT -16.690 139.250 -16.010 145.660 ;
        RECT -14.060 145.620 -13.590 145.660 ;
        RECT -11.890 142.460 -11.540 143.000 ;
        RECT 8.780 142.490 9.010 142.950 ;
        RECT -11.380 142.210 8.620 142.440 ;
        RECT -14.120 139.250 -13.680 139.360 ;
        RECT -16.690 138.710 -13.680 139.250 ;
        RECT -16.670 138.520 -13.680 138.710 ;
        RECT -14.120 138.390 -13.680 138.520 ;
        RECT -11.960 138.400 -11.470 139.390 ;
        RECT -11.840 137.100 -11.550 138.400 ;
        RECT -11.320 137.360 -10.760 142.210 ;
        RECT -3.680 137.360 -2.740 142.210 ;
        RECT 7.690 139.110 8.550 142.210 ;
        RECT 14.080 139.110 14.710 139.150 ;
        RECT 7.690 139.070 17.380 139.110 ;
        RECT 7.690 138.510 17.430 139.070 ;
        RECT 7.690 137.360 8.550 138.510 ;
        RECT -11.380 137.130 8.620 137.360 ;
        RECT -11.880 136.600 -11.540 137.100 ;
        RECT 8.780 136.620 9.010 137.080 ;
        RECT -11.840 136.550 -11.550 136.600 ;
        RECT 14.080 134.660 14.710 138.510 ;
        RECT 16.810 137.090 17.430 138.510 ;
        RECT 16.100 136.250 16.480 136.930 ;
        RECT 16.635 136.860 36.635 137.090 ;
        RECT 36.840 136.350 37.070 136.810 ;
        RECT 14.080 133.950 16.510 134.660 ;
        RECT 14.080 133.310 14.710 133.950 ;
        RECT 13.850 132.240 15.090 133.310 ;
        RECT -11.930 130.280 -11.570 130.800 ;
        RECT 8.730 130.320 8.960 130.780 ;
        RECT -11.430 130.040 8.570 130.270 ;
        RECT 16.050 130.080 16.510 133.950 ;
        RECT 36.900 130.160 37.130 130.620 ;
        RECT -3.680 125.240 -2.740 130.040 ;
        RECT 7.690 127.950 8.310 130.040 ;
        RECT 16.695 129.880 36.695 130.110 ;
        RECT 16.850 127.950 17.360 129.880 ;
        RECT 7.690 127.030 17.360 127.950 ;
        RECT 7.690 125.240 8.310 127.030 ;
        RECT -11.640 125.010 8.360 125.240 ;
        RECT -17.660 124.960 -11.830 124.990 ;
        RECT -17.660 124.510 -11.800 124.960 ;
        RECT -17.650 124.500 -11.800 124.510 ;
        RECT 8.520 124.500 8.750 124.960 ;
        RECT -17.650 124.420 -11.810 124.500 ;
        RECT 15.580 122.250 16.210 127.030 ;
        RECT 60.270 124.560 60.880 151.060 ;
        RECT 74.710 150.810 74.960 151.070 ;
        RECT 73.190 150.790 73.330 150.800 ;
        RECT 74.460 150.790 74.960 150.810 ;
        RECT 73.190 150.760 76.230 150.790 ;
        RECT 73.190 150.560 76.240 150.760 ;
        RECT 73.210 150.370 76.240 150.560 ;
        RECT 71.680 149.000 71.920 149.390 ;
        RECT 73.210 149.340 73.450 150.370 ;
        RECT 72.070 148.860 73.070 149.090 ;
        RECT 73.210 149.050 73.460 149.340 ;
        RECT 73.210 148.960 73.450 149.050 ;
        RECT 72.080 148.760 73.070 148.860 ;
        RECT 61.240 145.820 61.920 145.860 ;
        RECT 63.870 145.820 64.340 145.880 ;
        RECT 61.240 145.230 64.340 145.820 ;
        RECT 74.460 145.750 74.740 150.370 ;
        RECT 75.980 148.940 76.240 150.370 ;
        RECT 77.650 149.300 77.850 149.340 ;
        RECT 76.420 149.050 77.460 149.060 ;
        RECT 76.415 148.820 77.460 149.050 ;
        RECT 77.620 149.010 77.850 149.300 ;
        RECT 77.650 148.950 77.850 149.010 ;
        RECT 76.420 148.730 77.460 148.820 ;
        RECT 76.460 148.720 77.460 148.730 ;
        RECT 66.310 145.270 74.740 145.750 ;
        RECT 66.310 145.260 74.470 145.270 ;
        RECT 66.400 145.250 74.440 145.260 ;
        RECT 61.240 138.820 61.920 145.230 ;
        RECT 63.870 145.190 64.340 145.230 ;
        RECT 66.040 142.030 66.390 142.570 ;
        RECT 86.710 142.060 86.940 142.520 ;
        RECT 66.550 141.780 86.550 142.010 ;
        RECT 63.810 138.820 64.250 138.930 ;
        RECT 61.240 138.280 64.250 138.820 ;
        RECT 61.260 138.090 64.250 138.280 ;
        RECT 63.810 137.960 64.250 138.090 ;
        RECT 65.970 137.970 66.460 138.960 ;
        RECT 66.090 136.670 66.380 137.970 ;
        RECT 66.610 136.930 67.170 141.780 ;
        RECT 74.250 136.930 75.190 141.780 ;
        RECT 85.620 138.680 86.480 141.780 ;
        RECT 92.010 138.680 92.640 138.720 ;
        RECT 85.620 138.640 95.310 138.680 ;
        RECT 85.620 138.080 95.360 138.640 ;
        RECT 85.620 136.930 86.480 138.080 ;
        RECT 66.550 136.700 86.550 136.930 ;
        RECT 66.050 136.170 66.390 136.670 ;
        RECT 86.710 136.190 86.940 136.650 ;
        RECT 66.090 136.120 66.380 136.170 ;
        RECT 92.010 134.230 92.640 138.080 ;
        RECT 94.740 136.660 95.360 138.080 ;
        RECT 94.030 135.820 94.410 136.500 ;
        RECT 94.565 136.430 114.565 136.660 ;
        RECT 114.770 135.920 115.000 136.380 ;
        RECT 92.010 133.520 94.440 134.230 ;
        RECT 92.010 132.880 92.640 133.520 ;
        RECT 91.780 131.810 93.020 132.880 ;
        RECT 66.000 129.850 66.360 130.370 ;
        RECT 86.660 129.890 86.890 130.350 ;
        RECT 66.500 129.610 86.500 129.840 ;
        RECT 93.980 129.650 94.440 133.520 ;
        RECT 114.830 129.730 115.060 130.190 ;
        RECT 74.250 124.810 75.190 129.610 ;
        RECT 85.620 127.520 86.240 129.610 ;
        RECT 94.625 129.450 114.625 129.680 ;
        RECT 94.780 127.520 95.290 129.450 ;
        RECT 85.620 126.600 95.290 127.520 ;
        RECT 85.620 124.810 86.240 126.600 ;
        RECT 66.290 124.580 86.290 124.810 ;
        RECT 60.270 124.530 66.100 124.560 ;
        RECT 60.270 124.080 66.130 124.530 ;
        RECT 60.280 124.070 66.130 124.080 ;
        RECT 86.450 124.070 86.680 124.530 ;
        RECT 60.280 123.990 66.120 124.070 ;
        RECT 15.260 121.180 16.500 122.250 ;
        RECT 93.510 121.820 94.140 126.600 ;
        RECT 93.190 120.750 94.430 121.820 ;
        RECT 13.580 114.740 14.900 116.960 ;
        RECT 13.970 106.290 14.860 114.740 ;
        RECT 17.960 114.030 19.410 116.670 ;
        RECT -3.160 106.200 15.370 106.290 ;
        RECT 18.370 106.220 18.970 114.030 ;
        RECT -3.170 105.590 15.370 106.200 ;
        RECT -9.410 86.550 -8.980 86.620 ;
        RECT -3.170 86.550 -2.810 105.590 ;
        RECT 13.970 105.430 14.860 105.590 ;
        RECT 17.890 104.400 19.640 106.220 ;
        RECT 63.490 87.750 63.980 87.960 ;
        RECT 63.490 87.230 65.240 87.750 ;
        RECT 85.650 87.240 85.880 87.700 ;
        RECT 63.490 86.910 63.980 87.230 ;
        RECT 65.445 86.960 85.445 87.190 ;
        RECT -9.410 86.460 -2.810 86.550 ;
        RECT -9.410 86.120 -1.320 86.460 ;
        RECT -9.410 69.350 -8.980 86.120 ;
        RECT -3.170 85.940 -1.320 86.120 ;
        RECT 19.090 85.950 19.320 86.410 ;
        RECT -3.170 85.800 -2.810 85.940 ;
        RECT -1.115 85.670 18.885 85.900 ;
        RECT 62.900 85.880 63.080 85.890 ;
        RECT 65.630 85.880 66.980 86.960 ;
        RECT -3.660 84.590 -3.480 84.600 ;
        RECT -0.930 84.590 0.420 85.670 ;
        RECT -3.660 83.840 0.420 84.590 ;
        RECT -3.660 81.240 -3.480 83.840 ;
        RECT -2.970 82.800 -2.360 83.270 ;
        RECT -0.930 83.040 0.420 83.840 ;
        RECT 62.900 85.130 66.980 85.880 ;
        RECT -1.310 82.810 18.690 83.040 ;
        RECT -2.970 82.280 -1.470 82.800 ;
        RECT 18.850 82.300 19.080 82.760 ;
        RECT 62.900 82.670 63.080 85.130 ;
        RECT 65.630 84.330 66.980 85.130 ;
        RECT 63.590 84.090 64.280 84.260 ;
        RECT 65.250 84.100 85.250 84.330 ;
        RECT 63.590 83.570 65.090 84.090 ;
        RECT 85.410 83.590 85.640 84.050 ;
        RECT 63.590 83.450 64.280 83.570 ;
        RECT -2.970 81.890 -2.360 82.280 ;
        RECT 62.320 82.090 63.080 82.670 ;
        RECT 62.320 81.840 63.030 82.090 ;
        RECT -9.460 55.520 -8.980 69.350 ;
        RECT -227.980 44.500 -227.660 44.550 ;
        RECT -227.980 44.490 -200.680 44.500 ;
        RECT -227.980 43.890 -200.590 44.490 ;
        RECT -227.980 41.590 -227.660 43.890 ;
        RECT -222.460 43.510 -214.880 43.530 ;
        RECT -222.460 42.850 -214.690 43.510 ;
        RECT -233.860 30.130 -233.020 30.170 ;
        RECT -227.970 30.130 -227.670 41.590 ;
        RECT -222.420 40.900 -221.830 42.850 ;
        RECT -215.420 40.960 -214.690 42.850 ;
        RECT -222.480 40.430 -221.790 40.900 ;
        RECT -215.530 40.520 -214.560 40.960 ;
        RECT -222.350 38.370 -221.860 38.460 ;
        RECT -219.170 38.380 -218.630 38.730 ;
        RECT -215.560 38.680 -214.570 38.800 ;
        RECT -213.270 38.680 -212.770 38.720 ;
        RECT -215.560 38.390 -212.720 38.680 ;
        RECT -206.970 38.410 -206.450 38.770 ;
        RECT -201.160 38.670 -200.590 43.890 ;
        RECT -9.460 40.350 -9.030 55.520 ;
        RECT -201.130 38.650 -200.590 38.670 ;
        RECT -201.130 38.640 -200.670 38.650 ;
        RECT -225.990 32.850 -225.600 33.090 ;
        RECT -225.690 32.690 -225.460 32.700 ;
        RECT -225.690 31.700 -225.360 32.690 ;
        RECT -227.400 31.560 -227.160 31.580 ;
        RECT -227.400 31.440 -225.560 31.560 ;
        RECT -227.390 31.320 -225.560 31.440 ;
        RECT -227.390 30.310 -226.970 31.320 ;
        RECT -225.940 31.310 -225.650 31.320 ;
        RECT -222.350 30.330 -221.850 38.370 ;
        RECT -215.560 38.310 -214.570 38.390 ;
        RECT -213.270 38.380 -212.770 38.390 ;
        RECT -218.610 38.160 -218.380 38.220 ;
        RECT -213.530 38.160 -213.300 38.220 ;
        RECT -218.610 37.600 -213.300 38.160 ;
        RECT -218.610 30.520 -218.380 37.600 ;
        RECT -213.530 30.520 -213.300 37.600 ;
        RECT -222.350 30.310 -221.860 30.330 ;
        RECT -233.860 30.060 -227.670 30.130 ;
        RECT -227.410 30.300 -221.860 30.310 ;
        RECT -227.410 30.060 -221.870 30.300 ;
        RECT -233.860 30.030 -221.870 30.060 ;
        RECT -233.860 29.810 -226.970 30.030 ;
        RECT -233.860 29.800 -227.940 29.810 ;
        RECT -242.330 -4.430 -238.290 -4.170 ;
        RECT -242.330 -6.240 -236.320 -4.430 ;
        RECT -233.860 -6.240 -233.020 29.800 ;
        RECT -227.390 28.790 -226.970 29.810 ;
        RECT -218.610 29.580 -213.300 30.520 ;
        RECT -227.390 28.540 -225.540 28.790 ;
        RECT -227.360 28.530 -225.540 28.540 ;
        RECT -225.650 28.350 -225.420 28.355 ;
        RECT -225.660 28.310 -225.330 28.350 ;
        RECT -225.660 27.310 -225.320 28.310 ;
        RECT -225.900 27.120 -225.610 27.150 ;
        RECT -225.940 26.920 -225.550 27.120 ;
        RECT -218.610 19.150 -218.380 29.580 ;
        RECT -213.530 19.150 -213.300 29.580 ;
        RECT -218.610 18.290 -213.300 19.150 ;
        RECT -218.610 18.220 -218.380 18.290 ;
        RECT -219.120 17.830 -218.660 18.060 ;
        RECT -215.280 12.760 -214.680 18.290 ;
        RECT -213.530 18.220 -213.300 18.290 ;
        RECT -206.440 30.520 -206.210 38.270 ;
        RECT -201.410 30.520 -201.180 38.480 ;
        RECT -10.100 38.100 -8.250 40.350 ;
        RECT -116.520 36.300 -114.270 36.940 ;
        RECT -145.520 36.250 -114.270 36.300 ;
        RECT -162.790 35.870 -114.270 36.250 ;
        RECT -162.790 35.820 -131.690 35.870 ;
        RECT -206.440 29.580 -201.180 30.520 ;
        RECT -162.720 30.010 -162.290 35.820 ;
        RECT -116.520 35.090 -114.270 35.870 ;
        RECT -3.700 32.720 -3.320 81.240 ;
        RECT 12.540 59.730 15.530 63.200 ;
        RECT 13.610 55.290 14.430 59.730 ;
        RECT 0.330 54.530 14.650 55.290 ;
        RECT 0.540 37.920 1.020 54.530 ;
        RECT 85.580 45.850 87.685 46.750 ;
        RECT 20.890 43.310 22.995 44.210 ;
        RECT 86.550 43.530 87.110 45.850 ;
        RECT 21.690 40.540 22.080 43.310 ;
        RECT 86.350 43.150 87.260 43.530 ;
        RECT 86.350 43.130 90.290 43.150 ;
        RECT 86.350 42.760 90.300 43.130 ;
        RECT 86.340 42.440 90.300 42.760 ;
        RECT 86.340 41.420 87.260 42.440 ;
        RECT 65.330 40.650 65.850 40.990 ;
        RECT 86.340 40.880 87.250 41.420 ;
        RECT 67.295 40.650 87.295 40.880 ;
        RECT 21.530 40.160 22.440 40.540 ;
        RECT 21.530 40.140 25.470 40.160 ;
        RECT 21.530 39.770 25.480 40.140 ;
        RECT 65.330 40.130 67.090 40.650 ;
        RECT 87.500 40.140 87.730 40.600 ;
        RECT 65.330 39.950 65.850 40.130 ;
        RECT 67.295 39.860 87.295 40.090 ;
        RECT 0.270 37.660 1.020 37.920 ;
        RECT 21.520 39.450 25.480 39.770 ;
        RECT 21.520 38.430 22.440 39.450 ;
        RECT 21.520 37.890 22.430 38.430 ;
        RECT 2.475 37.660 22.475 37.890 ;
        RECT 0.270 37.140 2.270 37.660 ;
        RECT 22.680 37.150 22.910 37.610 ;
        RECT 0.270 36.930 0.890 37.140 ;
        RECT 2.475 36.870 22.475 37.100 ;
        RECT -0.070 35.790 0.110 35.800 ;
        RECT 2.660 35.790 4.010 36.870 ;
        RECT -0.070 35.040 4.010 35.790 ;
        RECT -4.330 32.160 -2.990 32.720 ;
        RECT -0.070 32.160 0.110 35.040 ;
        RECT 2.660 34.240 4.010 35.040 ;
        RECT 0.610 34.000 1.030 34.140 ;
        RECT 2.280 34.010 22.280 34.240 ;
        RECT 0.610 33.480 2.120 34.000 ;
        RECT 22.440 33.500 22.670 33.960 ;
        RECT 0.610 33.240 1.030 33.480 ;
        RECT 2.280 33.220 22.280 33.450 ;
        RECT 21.840 32.160 22.190 33.220 ;
        RECT 24.790 32.160 25.480 39.450 ;
        RECT 64.190 38.780 65.220 39.110 ;
        RECT 67.480 38.780 68.830 39.860 ;
        RECT 64.190 38.030 68.830 38.780 ;
        RECT 64.190 37.420 65.220 38.030 ;
        RECT 64.550 36.060 64.930 37.420 ;
        RECT 67.480 37.230 68.830 38.030 ;
        RECT 65.390 36.990 65.890 37.130 ;
        RECT 67.100 37.000 87.100 37.230 ;
        RECT 65.390 36.470 66.940 36.990 ;
        RECT 87.260 36.490 87.490 36.950 ;
        RECT 65.390 36.240 65.890 36.470 ;
        RECT 67.100 36.210 87.100 36.440 ;
        RECT 63.610 33.680 65.180 36.060 ;
        RECT 86.660 35.150 87.010 36.210 ;
        RECT 89.610 35.150 90.300 42.440 ;
        RECT 86.550 34.300 90.300 35.150 ;
        RECT 86.550 34.290 90.180 34.300 ;
        RECT -4.330 32.000 0.110 32.160 ;
        RECT -4.330 31.900 0.070 32.000 ;
        RECT -4.330 31.190 -2.990 31.900 ;
        RECT 21.730 31.310 25.480 32.160 ;
        RECT 21.730 31.300 25.360 31.310 ;
        RECT -108.890 30.540 -107.360 31.170 ;
        RECT -157.410 30.500 -107.360 30.540 ;
        RECT -160.770 30.320 -107.360 30.500 ;
        RECT -182.370 30.000 -161.970 30.010 ;
        RECT -206.440 19.150 -206.210 29.580 ;
        RECT -201.410 19.150 -201.180 29.580 ;
        RECT -206.440 18.530 -201.180 19.150 ;
        RECT -206.440 18.270 -206.210 18.530 ;
        RECT -213.250 17.830 -212.790 18.060 ;
        RECT -206.950 17.880 -206.490 18.110 ;
        RECT -209.480 12.760 -208.410 12.990 ;
        RECT -215.320 12.130 -208.410 12.760 ;
        RECT -215.280 10.030 -214.680 12.130 ;
        RECT -210.830 10.790 -210.120 12.130 ;
        RECT -209.480 11.750 -208.410 12.130 ;
        RECT -204.120 11.260 -203.200 18.530 ;
        RECT -201.410 18.480 -201.180 18.530 ;
        RECT -182.460 29.650 -161.970 30.000 ;
        RECT -201.130 18.090 -200.670 18.320 ;
        RECT -193.130 12.870 -190.910 13.260 ;
        RECT -182.460 12.870 -181.760 29.650 ;
        RECT -162.630 28.160 -162.110 29.650 ;
        RECT -162.070 27.770 -161.840 27.955 ;
        RECT -160.760 27.770 -160.010 30.320 ;
        RECT -157.410 30.160 -107.360 30.320 ;
        RECT -108.890 29.830 -107.360 30.160 ;
        RECT -159.440 29.200 -158.060 29.810 ;
        RECT -158.970 28.310 -158.450 29.200 ;
        RECT -159.210 27.770 -158.980 28.150 ;
        RECT -162.070 26.420 -158.980 27.770 ;
        RECT -108.330 26.910 -108.070 29.830 ;
        RECT 64.010 29.700 64.640 33.680 ;
        RECT 63.280 27.480 65.080 29.700 ;
        RECT -111.970 26.770 -108.070 26.910 ;
        RECT -111.970 26.730 -108.170 26.770 ;
        RECT -193.130 11.980 -181.600 12.870 ;
        RECT -193.130 11.940 -190.910 11.980 ;
        RECT -198.420 11.260 -197.350 11.580 ;
        RECT -182.460 11.470 -181.760 11.980 ;
        RECT -213.100 10.360 -212.420 10.740 ;
        RECT -210.830 10.330 -206.250 10.790 ;
        RECT -204.120 10.630 -197.350 11.260 ;
        RECT -213.260 10.030 -213.030 10.205 ;
        RECT -215.280 9.460 -213.030 10.030 ;
        RECT -215.240 9.410 -213.030 9.460 ;
        RECT -242.330 -6.700 -233.020 -6.240 ;
        RECT -242.330 -7.240 -238.290 -6.700 ;
        RECT -236.960 -6.870 -233.020 -6.700 ;
        RECT -233.860 -6.900 -233.020 -6.870 ;
        RECT -213.260 -9.795 -213.030 9.410 ;
        RECT -206.280 9.990 -206.050 10.145 ;
        RECT -204.120 9.990 -203.200 10.630 ;
        RECT -198.420 10.340 -197.350 10.630 ;
        RECT -206.280 9.480 -203.200 9.990 ;
        RECT -206.280 -9.855 -206.050 9.480 ;
        RECT -192.840 8.470 -190.200 8.880 ;
        RECT -182.390 8.470 -180.570 8.950 ;
        RECT -192.840 7.870 -180.570 8.470 ;
        RECT -162.070 7.955 -161.840 26.420 ;
        RECT -159.210 8.150 -158.980 26.420 ;
        RECT -131.460 26.300 -130.700 26.510 ;
        RECT -114.090 26.300 -113.100 26.570 ;
        RECT -131.460 25.950 -113.100 26.300 ;
        RECT -131.460 25.820 -113.310 25.950 ;
        RECT -139.370 13.230 -135.900 14.300 ;
        RECT -131.460 13.230 -130.700 25.820 ;
        RECT -113.830 24.570 -113.310 25.820 ;
        RECT -139.370 12.410 -130.700 13.230 ;
        RECT -139.370 11.310 -135.900 12.410 ;
        RECT -131.460 12.190 -130.700 12.410 ;
        RECT -192.840 7.430 -190.200 7.870 ;
        RECT -182.390 7.200 -180.570 7.870 ;
        RECT -158.930 7.760 -158.470 7.990 ;
        RECT -162.580 7.520 -162.120 7.750 ;
        RECT -120.380 5.150 -119.480 5.950 ;
        RECT -114.060 5.320 -113.830 24.365 ;
        RECT -115.940 5.310 -113.830 5.320 ;
        RECT -116.710 5.150 -113.830 5.310 ;
        RECT -120.380 4.760 -113.830 5.150 ;
        RECT -120.380 3.845 -119.480 4.760 ;
        RECT -116.710 4.410 -113.830 4.760 ;
        RECT -116.710 4.400 -114.600 4.410 ;
        RECT -116.330 2.050 -115.620 4.400 ;
        RECT -114.060 4.365 -113.830 4.410 ;
        RECT -113.270 24.180 -113.040 24.365 ;
        RECT -111.960 24.180 -111.210 26.730 ;
        RECT -110.310 25.810 -109.410 26.230 ;
        RECT -110.170 24.720 -109.650 25.810 ;
        RECT -110.410 24.180 -110.180 24.560 ;
        RECT -113.270 22.830 -110.180 24.180 ;
        RECT -113.270 4.365 -113.040 22.830 ;
        RECT -110.410 4.560 -110.180 22.830 ;
        RECT -109.620 5.000 -109.390 24.560 ;
        RECT -10.590 6.810 -9.900 6.960 ;
        RECT -10.670 6.750 0.340 6.810 ;
        RECT -10.670 6.660 6.415 6.750 ;
        RECT -10.670 6.470 6.420 6.660 ;
        RECT -10.670 6.340 2.340 6.470 ;
        RECT 4.120 6.360 6.420 6.470 ;
        RECT -10.670 6.270 0.340 6.340 ;
        RECT -108.330 5.000 -107.470 5.110 ;
        RECT -109.620 4.650 -107.470 5.000 ;
        RECT -109.620 4.560 -109.390 4.650 ;
        RECT -110.130 4.170 -109.670 4.400 ;
        RECT -113.780 3.930 -113.320 4.160 ;
        RECT -108.330 2.050 -107.470 4.650 ;
        RECT -116.330 1.480 -107.470 2.050 ;
        RECT -116.330 1.370 -107.480 1.480 ;
        RECT -116.310 1.360 -107.480 1.370 ;
        RECT -10.590 -7.270 -9.900 6.270 ;
        RECT 1.740 4.440 2.340 6.340 ;
        RECT 3.340 4.440 3.940 6.240 ;
        RECT 5.820 4.460 6.420 6.360 ;
        RECT 7.420 4.460 8.020 6.260 ;
        RECT -1.550 4.110 -0.840 4.240 ;
        RECT 2.340 4.140 3.340 4.240 ;
        RECT 6.420 4.160 7.420 4.260 ;
        RECT 4.220 4.140 8.020 4.160 ;
        RECT 0.135 4.110 8.020 4.140 ;
        RECT -1.550 3.860 8.020 4.110 ;
        RECT -1.550 3.840 3.940 3.860 ;
        RECT -1.550 3.790 0.400 3.840 ;
        RECT -1.550 3.600 -0.840 3.790 ;
        RECT -5.090 3.260 -4.580 3.280 ;
        RECT -5.090 3.200 0.430 3.260 ;
        RECT 4.060 3.200 6.360 3.220 ;
        RECT -5.090 2.955 6.360 3.200 ;
        RECT -5.090 2.900 2.300 2.955 ;
        RECT 4.060 2.920 6.360 2.955 ;
        RECT -5.090 2.890 0.430 2.900 ;
        RECT -5.090 -1.200 -4.580 2.890 ;
        RECT 1.700 1.000 2.300 2.900 ;
        RECT 3.300 1.000 3.900 2.800 ;
        RECT 5.760 1.020 6.360 2.920 ;
        RECT 7.360 1.020 7.960 2.820 ;
        RECT -1.630 0.700 -0.920 0.890 ;
        RECT 2.300 0.700 3.300 0.800 ;
        RECT 6.360 0.720 7.360 0.820 ;
        RECT 4.160 0.700 7.960 0.720 ;
        RECT -1.630 0.420 7.960 0.700 ;
        RECT -1.630 0.400 3.900 0.420 ;
        RECT -1.630 0.380 0.320 0.400 ;
        RECT -1.630 0.250 -0.920 0.380 ;
        RECT 63.440 -1.190 66.990 -1.040 ;
        RECT 5.820 -1.200 66.990 -1.190 ;
        RECT -5.090 -1.720 66.990 -1.200 ;
        RECT -5.050 -1.740 66.990 -1.720 ;
        RECT 5.820 -1.780 66.990 -1.740 ;
        RECT 63.440 -2.060 66.990 -1.780 ;
        RECT -1.770 -7.270 -0.970 -7.240 ;
        RECT -10.590 -8.000 -0.950 -7.270 ;
        RECT -10.430 -8.040 -0.950 -8.000 ;
        RECT -212.980 -10.230 -212.520 -10.000 ;
        RECT -206.790 -10.290 -206.330 -10.060 ;
        RECT -287.110 -15.970 -286.880 -15.340 ;
        RECT -279.910 -15.950 -278.200 -15.940 ;
        RECT -275.990 -15.950 -275.660 -15.910 ;
        RECT -287.110 -16.240 -285.260 -15.970 ;
        RECT -287.110 -16.340 -286.880 -16.240 ;
        RECT -285.490 -17.660 -285.260 -16.240 ;
        RECT -279.910 -16.190 -275.660 -15.950 ;
        RECT -267.620 -16.080 -267.290 -15.800 ;
        RECT -285.490 -17.940 -280.710 -17.660 ;
        RECT -287.060 -18.980 -286.830 -18.705 ;
        RECT -285.490 -18.980 -285.260 -17.940 ;
        RECT -281.150 -18.330 -280.710 -17.940 ;
        RECT -279.910 -18.330 -279.360 -16.190 ;
        RECT -278.700 -16.200 -275.660 -16.190 ;
        RECT -275.970 -16.210 -275.680 -16.200 ;
        RECT -247.330 -16.240 -247.000 -15.960 ;
        RECT -276.160 -16.980 -275.930 -16.370 ;
        RECT -277.440 -17.240 -275.930 -16.980 ;
        RECT -281.150 -18.880 -279.360 -18.330 ;
        RECT -277.430 -18.480 -277.070 -17.240 ;
        RECT -276.160 -17.370 -275.930 -17.240 ;
        RECT -275.720 -16.810 -275.490 -16.370 ;
        RECT -272.700 -16.810 -272.470 -16.260 ;
        RECT -275.720 -17.100 -272.470 -16.810 ;
        RECT -275.720 -17.370 -275.490 -17.100 ;
        RECT -272.700 -17.260 -272.470 -17.100 ;
        RECT -267.350 -16.790 -267.120 -16.240 ;
        RECT -267.350 -16.830 -265.470 -16.790 ;
        RECT -267.350 -17.120 -265.390 -16.830 ;
        RECT -267.350 -17.240 -267.120 -17.120 ;
        RECT -275.990 -17.800 -275.660 -17.520 ;
        RECT -267.710 -17.770 -267.150 -17.390 ;
        RECT -265.620 -18.410 -265.390 -17.120 ;
        RECT -255.870 -17.140 -255.640 -16.530 ;
        RECT -257.150 -17.400 -255.640 -17.140 ;
        RECT -278.230 -18.520 -272.860 -18.480 ;
        RECT -278.230 -18.750 -270.860 -18.520 ;
        RECT -281.150 -18.900 -280.710 -18.880 ;
        RECT -287.060 -19.240 -285.260 -18.980 ;
        RECT -287.060 -19.705 -286.830 -19.240 ;
        RECT -279.910 -21.270 -279.360 -18.880 ;
        RECT -278.190 -20.200 -277.920 -18.750 ;
        RECT -276.230 -18.790 -270.860 -18.750 ;
        RECT -274.550 -19.300 -273.610 -18.790 ;
        RECT -275.960 -19.840 -275.630 -19.560 ;
        RECT -275.950 -19.850 -275.660 -19.840 ;
        RECT -276.140 -20.200 -275.910 -20.055 ;
        RECT -278.190 -20.320 -275.910 -20.200 ;
        RECT -278.160 -20.340 -275.910 -20.320 ;
        RECT -276.140 -21.055 -275.910 -20.340 ;
        RECT -272.280 -20.260 -272.050 -20.075 ;
        RECT -271.170 -20.260 -270.870 -18.790 ;
        RECT -267.660 -19.950 -267.160 -19.610 ;
        RECT -265.620 -19.650 -263.980 -18.410 ;
        RECT -257.140 -18.640 -256.780 -17.400 ;
        RECT -255.870 -17.530 -255.640 -17.400 ;
        RECT -255.430 -16.970 -255.200 -16.530 ;
        RECT -252.410 -16.970 -252.180 -16.420 ;
        RECT -255.430 -17.260 -252.180 -16.970 ;
        RECT -255.430 -17.530 -255.200 -17.260 ;
        RECT -252.410 -17.420 -252.180 -17.260 ;
        RECT -247.060 -16.950 -246.830 -16.400 ;
        RECT -247.060 -16.990 -245.180 -16.950 ;
        RECT -247.060 -17.280 -245.100 -16.990 ;
        RECT -247.060 -17.400 -246.830 -17.280 ;
        RECT -247.420 -17.930 -246.860 -17.550 ;
        RECT -245.330 -18.040 -245.100 -17.280 ;
        RECT -257.940 -18.680 -252.570 -18.640 ;
        RECT -257.940 -18.910 -250.570 -18.680 ;
        RECT -272.280 -20.480 -270.870 -20.260 ;
        RECT -267.290 -20.170 -267.060 -20.145 ;
        RECT -265.620 -20.170 -265.390 -19.650 ;
        RECT -272.280 -21.075 -272.050 -20.480 ;
        RECT -267.290 -20.500 -265.390 -20.170 ;
        RECT -257.900 -20.360 -257.630 -18.910 ;
        RECT -255.940 -18.950 -250.570 -18.910 ;
        RECT -254.260 -19.460 -253.320 -18.950 ;
        RECT -255.850 -20.360 -255.620 -20.215 ;
        RECT -257.900 -20.480 -255.620 -20.360 ;
        RECT -257.870 -20.500 -255.620 -20.480 ;
        RECT -267.290 -21.145 -267.060 -20.500 ;
        RECT -255.850 -21.215 -255.620 -20.500 ;
        RECT -251.990 -20.420 -251.760 -20.235 ;
        RECT -250.880 -20.420 -250.580 -18.950 ;
        RECT -245.330 -19.450 -238.700 -18.040 ;
        RECT -247.370 -20.110 -246.870 -19.770 ;
        RECT -251.990 -20.640 -250.580 -20.420 ;
        RECT -247.000 -20.330 -246.770 -20.305 ;
        RECT -245.330 -20.330 -245.100 -19.450 ;
        RECT -251.990 -21.235 -251.760 -20.640 ;
        RECT -247.000 -20.660 -245.100 -20.330 ;
        RECT -275.960 -21.270 -275.630 -21.240 ;
        RECT -279.910 -21.580 -275.620 -21.270 ;
        RECT -247.000 -21.305 -246.770 -20.660 ;
        RECT -279.910 -21.590 -279.360 -21.580 ;
        RECT -267.560 -21.620 -267.230 -21.340 ;
        RECT -247.270 -21.780 -246.940 -21.500 ;
        RECT -239.590 -47.890 -238.760 -19.450 ;
        RECT -227.550 -33.430 -227.230 -33.380 ;
        RECT -227.550 -33.440 -200.250 -33.430 ;
        RECT -227.550 -34.040 -200.160 -33.440 ;
        RECT -227.550 -36.340 -227.230 -34.040 ;
        RECT -222.030 -34.420 -214.450 -34.400 ;
        RECT -222.030 -35.080 -214.260 -34.420 ;
        RECT -227.540 -47.870 -227.240 -36.340 ;
        RECT -221.990 -37.030 -221.400 -35.080 ;
        RECT -214.990 -36.970 -214.260 -35.080 ;
        RECT -222.050 -37.500 -221.360 -37.030 ;
        RECT -215.100 -37.410 -214.130 -36.970 ;
        RECT -221.920 -39.560 -221.430 -39.470 ;
        RECT -218.740 -39.550 -218.200 -39.200 ;
        RECT -215.130 -39.250 -214.140 -39.130 ;
        RECT -212.840 -39.250 -212.340 -39.210 ;
        RECT -215.130 -39.540 -212.290 -39.250 ;
        RECT -206.540 -39.520 -206.020 -39.160 ;
        RECT -200.730 -39.260 -200.160 -34.040 ;
        RECT -158.840 -36.060 -158.010 -35.480 ;
        RECT -162.060 -36.190 -158.010 -36.060 ;
        RECT -162.060 -36.240 -158.260 -36.190 ;
        RECT -164.130 -37.140 -163.080 -36.650 ;
        RECT -163.920 -38.400 -163.400 -37.140 ;
        RECT -200.700 -39.280 -200.160 -39.260 ;
        RECT -163.360 -38.790 -163.130 -38.605 ;
        RECT -162.050 -38.790 -161.300 -36.240 ;
        RECT -160.430 -37.440 -159.620 -36.750 ;
        RECT -112.230 -37.170 -109.850 -36.770 ;
        RECT -105.870 -37.170 -103.650 -36.440 ;
        RECT -160.260 -38.250 -159.740 -37.440 ;
        RECT -115.280 -37.710 -113.590 -37.350 ;
        RECT -112.230 -37.710 -103.650 -37.170 ;
        RECT -115.280 -37.800 -103.650 -37.710 ;
        RECT -115.280 -38.090 -109.850 -37.800 ;
        RECT -115.280 -38.380 -113.590 -38.090 ;
        RECT -112.230 -38.340 -109.850 -38.090 ;
        RECT -105.870 -38.240 -103.650 -37.800 ;
        RECT -160.500 -38.790 -160.270 -38.410 ;
        RECT -200.700 -39.290 -200.240 -39.280 ;
        RECT -225.560 -45.080 -225.170 -44.840 ;
        RECT -225.260 -45.240 -225.030 -45.230 ;
        RECT -225.260 -46.230 -224.930 -45.240 ;
        RECT -226.970 -46.370 -226.730 -46.350 ;
        RECT -226.970 -46.490 -225.130 -46.370 ;
        RECT -226.960 -46.610 -225.130 -46.490 ;
        RECT -226.960 -47.620 -226.540 -46.610 ;
        RECT -225.510 -46.620 -225.220 -46.610 ;
        RECT -221.920 -47.600 -221.420 -39.560 ;
        RECT -215.130 -39.620 -214.140 -39.540 ;
        RECT -212.840 -39.550 -212.340 -39.540 ;
        RECT -218.180 -39.770 -217.950 -39.710 ;
        RECT -213.100 -39.770 -212.870 -39.710 ;
        RECT -218.180 -40.330 -212.870 -39.770 ;
        RECT -218.180 -47.410 -217.950 -40.330 ;
        RECT -213.100 -47.410 -212.870 -40.330 ;
        RECT -221.920 -47.620 -221.430 -47.600 ;
        RECT -226.980 -47.630 -221.430 -47.620 ;
        RECT -226.980 -47.870 -221.440 -47.630 ;
        RECT -227.720 -47.890 -221.440 -47.870 ;
        RECT -239.590 -47.900 -221.440 -47.890 ;
        RECT -239.590 -48.120 -226.540 -47.900 ;
        RECT -239.590 -48.170 -227.600 -48.120 ;
        RECT -239.450 -48.180 -227.600 -48.170 ;
        RECT -226.960 -49.140 -226.540 -48.120 ;
        RECT -218.180 -48.350 -212.870 -47.410 ;
        RECT -226.960 -49.390 -225.110 -49.140 ;
        RECT -226.930 -49.400 -225.110 -49.390 ;
        RECT -225.220 -49.580 -224.990 -49.575 ;
        RECT -225.230 -49.620 -224.900 -49.580 ;
        RECT -225.230 -50.620 -224.890 -49.620 ;
        RECT -225.470 -50.810 -225.180 -50.780 ;
        RECT -225.510 -51.010 -225.120 -50.810 ;
        RECT -218.180 -58.780 -217.950 -48.350 ;
        RECT -213.100 -58.780 -212.870 -48.350 ;
        RECT -218.180 -59.640 -212.870 -58.780 ;
        RECT -218.180 -59.710 -217.950 -59.640 ;
        RECT -218.690 -60.100 -218.230 -59.870 ;
        RECT -214.850 -65.170 -214.250 -59.640 ;
        RECT -213.100 -59.710 -212.870 -59.640 ;
        RECT -206.010 -47.410 -205.780 -39.660 ;
        RECT -200.980 -47.410 -200.750 -39.450 ;
        RECT -206.010 -48.350 -200.750 -47.410 ;
        RECT -206.010 -58.780 -205.780 -48.350 ;
        RECT -200.980 -58.780 -200.750 -48.350 ;
        RECT -163.360 -40.140 -160.270 -38.790 ;
        RECT -117.160 -39.010 -116.120 -38.490 ;
        RECT -163.360 -58.605 -163.130 -40.140 ;
        RECT -160.500 -58.410 -160.270 -40.140 ;
        RECT -116.820 -40.250 -116.300 -39.010 ;
        RECT -206.010 -59.400 -200.750 -58.780 ;
        RECT -160.220 -58.800 -159.760 -58.570 ;
        RECT -163.870 -59.040 -163.410 -58.810 ;
        RECT -206.010 -59.660 -205.780 -59.400 ;
        RECT -212.820 -60.100 -212.360 -59.870 ;
        RECT -206.520 -60.050 -206.060 -59.820 ;
        RECT -209.050 -65.170 -207.980 -64.940 ;
        RECT -214.890 -65.800 -207.980 -65.170 ;
        RECT -214.850 -67.900 -214.250 -65.800 ;
        RECT -210.400 -67.140 -209.690 -65.800 ;
        RECT -209.050 -66.180 -207.980 -65.800 ;
        RECT -203.690 -66.670 -202.770 -59.400 ;
        RECT -200.980 -59.450 -200.750 -59.400 ;
        RECT -200.700 -59.840 -200.240 -59.610 ;
        RECT -122.920 -59.710 -122.020 -58.740 ;
        RECT -117.050 -59.500 -116.820 -40.455 ;
        RECT -118.930 -59.510 -116.820 -59.500 ;
        RECT -119.700 -59.710 -116.820 -59.510 ;
        RECT -122.920 -60.270 -116.820 -59.710 ;
        RECT -122.920 -60.845 -122.020 -60.270 ;
        RECT -119.700 -60.410 -116.820 -60.270 ;
        RECT -119.700 -60.420 -117.590 -60.410 ;
        RECT -119.320 -62.770 -118.610 -60.420 ;
        RECT -117.050 -60.455 -116.820 -60.410 ;
        RECT -116.260 -40.640 -116.030 -40.455 ;
        RECT -114.950 -40.640 -114.200 -38.380 ;
        RECT -113.300 -39.050 -112.410 -38.550 ;
        RECT -113.160 -40.100 -112.640 -39.050 ;
        RECT -113.400 -40.640 -113.170 -40.260 ;
        RECT -116.260 -41.990 -113.170 -40.640 ;
        RECT -116.260 -60.455 -116.030 -41.990 ;
        RECT -113.400 -60.260 -113.170 -41.990 ;
        RECT -112.610 -59.820 -112.380 -40.260 ;
        RECT -1.770 -44.520 -0.970 -8.040 ;
        RECT -2.050 -45.580 -0.670 -44.520 ;
        RECT 66.320 -45.310 66.960 -2.060 ;
        RECT 66.140 -45.930 67.070 -45.310 ;
        RECT 65.700 -55.590 67.500 -53.370 ;
        RECT -1.910 -57.790 -0.570 -57.080 ;
        RECT 24.150 -57.200 27.780 -57.190 ;
        RECT -1.910 -57.890 2.490 -57.790 ;
        RECT -1.910 -58.050 2.530 -57.890 ;
        RECT 24.150 -58.050 27.900 -57.200 ;
        RECT -1.910 -58.610 -0.570 -58.050 ;
        RECT -111.320 -59.820 -110.460 -59.710 ;
        RECT -112.610 -60.170 -110.460 -59.820 ;
        RECT -112.610 -60.260 -112.380 -60.170 ;
        RECT -113.120 -60.650 -112.660 -60.420 ;
        RECT -116.770 -60.890 -116.310 -60.660 ;
        RECT -111.320 -62.770 -110.460 -60.170 ;
        RECT -119.320 -63.340 -110.460 -62.770 ;
        RECT -119.320 -63.450 -110.470 -63.340 ;
        RECT -119.300 -63.460 -110.470 -63.450 ;
        RECT -7.680 -66.240 -5.830 -63.990 ;
        RECT -197.990 -66.670 -196.920 -66.350 ;
        RECT -212.670 -67.570 -211.990 -67.190 ;
        RECT -210.400 -67.600 -205.820 -67.140 ;
        RECT -203.690 -67.300 -196.920 -66.670 ;
        RECT -212.830 -67.900 -212.600 -67.725 ;
        RECT -214.850 -68.470 -212.600 -67.900 ;
        RECT -214.810 -68.520 -212.600 -68.470 ;
        RECT -212.830 -87.725 -212.600 -68.520 ;
        RECT -205.850 -67.940 -205.620 -67.785 ;
        RECT -203.690 -67.940 -202.770 -67.300 ;
        RECT -197.990 -67.590 -196.920 -67.300 ;
        RECT -205.850 -68.450 -202.770 -67.940 ;
        RECT -205.850 -87.785 -205.620 -68.450 ;
        RECT -7.040 -81.410 -6.610 -66.240 ;
        RECT -212.550 -88.160 -212.090 -87.930 ;
        RECT -206.360 -88.220 -205.900 -87.990 ;
        RECT -7.040 -95.240 -6.560 -81.410 ;
        RECT -6.990 -112.010 -6.560 -95.240 ;
        RECT -1.280 -107.130 -0.900 -58.610 ;
        RECT 2.350 -60.930 2.530 -58.050 ;
        RECT 24.260 -59.110 24.610 -58.050 ;
        RECT 3.030 -59.370 3.450 -59.130 ;
        RECT 4.700 -59.340 24.700 -59.110 ;
        RECT 3.030 -59.890 4.540 -59.370 ;
        RECT 24.860 -59.850 25.090 -59.390 ;
        RECT 3.030 -60.030 3.450 -59.890 ;
        RECT 4.700 -60.130 24.700 -59.900 ;
        RECT 5.080 -60.930 6.430 -60.130 ;
        RECT 2.350 -61.680 6.430 -60.930 ;
        RECT 2.350 -61.690 2.530 -61.680 ;
        RECT 5.080 -62.760 6.430 -61.680 ;
        RECT 2.690 -63.030 3.310 -62.820 ;
        RECT 4.895 -62.990 24.895 -62.760 ;
        RECT 2.690 -63.550 4.690 -63.030 ;
        RECT 25.100 -63.500 25.330 -63.040 ;
        RECT 2.690 -63.810 3.440 -63.550 ;
        RECT 4.895 -63.780 24.895 -63.550 ;
        RECT 2.960 -80.420 3.440 -63.810 ;
        RECT 23.940 -64.320 24.850 -63.780 ;
        RECT 23.940 -65.340 24.860 -64.320 ;
        RECT 27.210 -65.340 27.900 -58.050 ;
        RECT 66.430 -59.570 67.060 -55.590 ;
        RECT 66.030 -61.950 67.600 -59.570 ;
        RECT 88.970 -60.190 92.600 -60.180 ;
        RECT 88.970 -61.040 92.720 -60.190 ;
        RECT 66.970 -63.310 67.350 -61.950 ;
        RECT 89.080 -62.100 89.430 -61.040 ;
        RECT 67.810 -62.360 68.310 -62.130 ;
        RECT 69.520 -62.330 89.520 -62.100 ;
        RECT 67.810 -62.880 69.360 -62.360 ;
        RECT 89.680 -62.840 89.910 -62.380 ;
        RECT 67.810 -63.020 68.310 -62.880 ;
        RECT 69.520 -63.120 89.520 -62.890 ;
        RECT 66.610 -63.920 67.640 -63.310 ;
        RECT 69.900 -63.920 71.250 -63.120 ;
        RECT 66.610 -64.670 71.250 -63.920 ;
        RECT 66.610 -65.000 67.640 -64.670 ;
        RECT 23.940 -65.660 27.900 -65.340 ;
        RECT 23.950 -66.030 27.900 -65.660 ;
        RECT 69.900 -65.750 71.250 -64.670 ;
        RECT 67.750 -66.020 68.270 -65.840 ;
        RECT 69.715 -65.980 89.715 -65.750 ;
        RECT 23.950 -66.050 27.890 -66.030 ;
        RECT 23.950 -66.430 24.860 -66.050 ;
        RECT 24.110 -69.200 24.500 -66.430 ;
        RECT 67.750 -66.540 69.510 -66.020 ;
        RECT 89.920 -66.490 90.150 -66.030 ;
        RECT 67.750 -66.880 68.270 -66.540 ;
        RECT 69.715 -66.770 89.715 -66.540 ;
        RECT 88.760 -67.310 89.670 -66.770 ;
        RECT 88.760 -68.330 89.680 -67.310 ;
        RECT 92.030 -68.330 92.720 -61.040 ;
        RECT 88.760 -68.650 92.720 -68.330 ;
        RECT 88.770 -69.020 92.720 -68.650 ;
        RECT 88.770 -69.040 92.710 -69.020 ;
        RECT 23.310 -70.100 25.415 -69.200 ;
        RECT 88.770 -69.420 89.680 -69.040 ;
        RECT 88.970 -71.740 89.530 -69.420 ;
        RECT 88.000 -72.640 90.105 -71.740 ;
        RECT 2.750 -81.180 17.070 -80.420 ;
        RECT 16.030 -85.620 16.850 -81.180 ;
        RECT 14.960 -89.090 17.950 -85.620 ;
        RECT -1.240 -109.730 -1.060 -107.130 ;
        RECT -0.550 -108.170 0.060 -107.780 ;
        RECT 64.740 -107.980 65.450 -107.730 ;
        RECT -0.550 -108.690 0.950 -108.170 ;
        RECT 21.270 -108.650 21.500 -108.190 ;
        RECT 64.740 -108.560 65.500 -107.980 ;
        RECT -0.550 -109.160 0.060 -108.690 ;
        RECT 1.110 -108.930 21.110 -108.700 ;
        RECT 1.490 -109.730 2.840 -108.930 ;
        RECT -1.240 -110.480 2.840 -109.730 ;
        RECT -1.240 -110.490 -1.060 -110.480 ;
        RECT 1.490 -111.560 2.840 -110.480 ;
        RECT 65.320 -111.020 65.500 -108.560 ;
        RECT 66.010 -109.460 66.700 -109.340 ;
        RECT 66.010 -109.980 67.510 -109.460 ;
        RECT 87.830 -109.940 88.060 -109.480 ;
        RECT 66.010 -110.150 66.700 -109.980 ;
        RECT 67.670 -110.220 87.670 -109.990 ;
        RECT 68.050 -111.020 69.400 -110.220 ;
        RECT -0.750 -111.830 -0.390 -111.690 ;
        RECT 1.305 -111.790 21.305 -111.560 ;
        RECT 65.320 -111.770 69.400 -111.020 ;
        RECT 65.320 -111.780 65.500 -111.770 ;
        RECT -0.750 -112.010 1.100 -111.830 ;
        RECT -6.990 -112.350 1.100 -112.010 ;
        RECT 21.510 -112.300 21.740 -111.840 ;
        RECT -6.990 -112.440 -0.390 -112.350 ;
        RECT -6.990 -112.510 -6.560 -112.440 ;
        RECT -0.750 -131.480 -0.390 -112.440 ;
        RECT 65.910 -113.120 66.400 -112.800 ;
        RECT 68.050 -112.850 69.400 -111.770 ;
        RECT 67.865 -113.080 87.865 -112.850 ;
        RECT 65.910 -113.640 67.660 -113.120 ;
        RECT 88.070 -113.590 88.300 -113.130 ;
        RECT 65.910 -113.850 66.400 -113.640 ;
        RECT 16.390 -131.480 17.280 -131.320 ;
        RECT -0.750 -132.090 17.790 -131.480 ;
        RECT -0.740 -132.180 17.790 -132.090 ;
        RECT 20.310 -132.110 22.060 -130.290 ;
        RECT 16.390 -140.630 17.280 -132.180 ;
        RECT 20.790 -139.920 21.390 -132.110 ;
        RECT 16.000 -142.850 17.320 -140.630 ;
        RECT 20.380 -142.560 21.830 -139.920 ;
        RECT 17.680 -148.140 18.920 -147.070 ;
        RECT 95.610 -147.710 96.850 -146.640 ;
        RECT -15.230 -150.390 -9.390 -150.310 ;
        RECT -15.230 -150.400 -9.380 -150.390 ;
        RECT -15.240 -150.850 -9.380 -150.400 ;
        RECT 10.940 -150.850 11.170 -150.390 ;
        RECT -15.240 -150.880 -9.410 -150.850 ;
        RECT -15.240 -177.380 -14.630 -150.880 ;
        RECT -9.220 -151.130 10.780 -150.900 ;
        RECT -1.260 -155.930 -0.320 -151.130 ;
        RECT 10.110 -152.920 10.730 -151.130 ;
        RECT 18.000 -152.920 18.630 -148.140 ;
        RECT 62.700 -149.960 68.540 -149.880 ;
        RECT 62.700 -149.970 68.550 -149.960 ;
        RECT 62.690 -150.420 68.550 -149.970 ;
        RECT 88.870 -150.420 89.100 -149.960 ;
        RECT 62.690 -150.450 68.520 -150.420 ;
        RECT 10.110 -153.840 19.780 -152.920 ;
        RECT 10.110 -155.930 10.730 -153.840 ;
        RECT 19.270 -155.770 19.780 -153.840 ;
        RECT -9.010 -156.160 10.990 -155.930 ;
        RECT -9.510 -156.690 -9.150 -156.170 ;
        RECT 11.150 -156.670 11.380 -156.210 ;
        RECT 16.270 -159.200 17.510 -158.130 ;
        RECT 16.500 -159.840 17.130 -159.200 ;
        RECT 18.470 -159.840 18.930 -155.970 ;
        RECT 19.115 -156.000 39.115 -155.770 ;
        RECT 39.320 -156.510 39.550 -156.050 ;
        RECT 16.500 -160.550 18.930 -159.840 ;
        RECT -9.420 -162.490 -9.130 -162.440 ;
        RECT -9.460 -162.990 -9.120 -162.490 ;
        RECT 11.200 -162.970 11.430 -162.510 ;
        RECT -11.700 -164.410 -11.260 -164.280 ;
        RECT -9.420 -164.290 -9.130 -162.990 ;
        RECT -8.960 -163.250 11.040 -163.020 ;
        RECT -14.250 -164.600 -11.260 -164.410 ;
        RECT -14.270 -165.140 -11.260 -164.600 ;
        RECT -14.270 -171.550 -13.590 -165.140 ;
        RECT -11.700 -165.250 -11.260 -165.140 ;
        RECT -9.540 -165.280 -9.050 -164.290 ;
        RECT -8.900 -168.100 -8.340 -163.250 ;
        RECT -1.260 -168.100 -0.320 -163.250 ;
        RECT 10.110 -164.400 10.970 -163.250 ;
        RECT 16.500 -164.400 17.130 -160.550 ;
        RECT 18.520 -162.820 18.900 -162.140 ;
        RECT 39.260 -162.700 39.490 -162.240 ;
        RECT 19.055 -162.980 39.055 -162.750 ;
        RECT 19.230 -164.400 19.850 -162.980 ;
        RECT 10.110 -164.960 19.850 -164.400 ;
        RECT 10.110 -165.000 19.800 -164.960 ;
        RECT 10.110 -168.100 10.970 -165.000 ;
        RECT 16.500 -165.040 17.130 -165.000 ;
        RECT -8.960 -168.330 11.040 -168.100 ;
        RECT -9.470 -168.890 -9.120 -168.350 ;
        RECT 11.200 -168.840 11.430 -168.380 ;
        RECT -11.640 -171.550 -11.170 -171.510 ;
        RECT -14.270 -172.140 -11.170 -171.550 ;
        RECT -9.110 -171.580 -1.070 -171.570 ;
        RECT -9.200 -171.590 -1.040 -171.580 ;
        RECT -9.200 -172.070 -0.770 -171.590 ;
        RECT -14.270 -172.180 -13.590 -172.140 ;
        RECT -11.640 -172.200 -11.170 -172.140 ;
        RECT -3.430 -175.180 -2.440 -175.080 ;
        RECT -3.830 -175.710 -3.590 -175.320 ;
        RECT -3.440 -175.410 -2.440 -175.180 ;
        RECT -2.300 -175.370 -2.060 -175.280 ;
        RECT -2.300 -175.660 -2.050 -175.370 ;
        RECT -2.300 -176.690 -2.060 -175.660 ;
        RECT -1.050 -176.690 -0.770 -172.070 ;
        RECT 0.950 -175.050 1.950 -175.040 ;
        RECT 0.910 -175.140 1.950 -175.050 ;
        RECT 0.470 -176.690 0.730 -175.260 ;
        RECT 0.905 -175.370 1.950 -175.140 ;
        RECT 2.140 -175.330 2.340 -175.270 ;
        RECT 0.910 -175.380 1.950 -175.370 ;
        RECT 2.110 -175.620 2.340 -175.330 ;
        RECT 2.140 -175.660 2.340 -175.620 ;
        RECT -2.300 -176.880 0.730 -176.690 ;
        RECT -2.320 -177.080 0.730 -176.880 ;
        RECT 62.690 -176.950 63.300 -150.450 ;
        RECT 68.710 -150.700 88.710 -150.470 ;
        RECT 76.670 -155.500 77.610 -150.700 ;
        RECT 88.040 -152.490 88.660 -150.700 ;
        RECT 95.930 -152.490 96.560 -147.710 ;
        RECT 88.040 -153.410 97.710 -152.490 ;
        RECT 88.040 -155.500 88.660 -153.410 ;
        RECT 97.200 -155.340 97.710 -153.410 ;
        RECT 68.920 -155.730 88.920 -155.500 ;
        RECT 68.420 -156.260 68.780 -155.740 ;
        RECT 89.080 -156.240 89.310 -155.780 ;
        RECT 94.200 -158.770 95.440 -157.700 ;
        RECT 94.430 -159.410 95.060 -158.770 ;
        RECT 96.400 -159.410 96.860 -155.540 ;
        RECT 97.045 -155.570 117.045 -155.340 ;
        RECT 117.250 -156.080 117.480 -155.620 ;
        RECT 94.430 -160.120 96.860 -159.410 ;
        RECT 68.510 -162.060 68.800 -162.010 ;
        RECT 68.470 -162.560 68.810 -162.060 ;
        RECT 89.130 -162.540 89.360 -162.080 ;
        RECT 66.230 -163.980 66.670 -163.850 ;
        RECT 68.510 -163.860 68.800 -162.560 ;
        RECT 68.970 -162.820 88.970 -162.590 ;
        RECT 63.680 -164.170 66.670 -163.980 ;
        RECT 63.660 -164.710 66.670 -164.170 ;
        RECT 63.660 -171.120 64.340 -164.710 ;
        RECT 66.230 -164.820 66.670 -164.710 ;
        RECT 68.390 -164.850 68.880 -163.860 ;
        RECT 69.030 -167.670 69.590 -162.820 ;
        RECT 76.670 -167.670 77.610 -162.820 ;
        RECT 88.040 -163.970 88.900 -162.820 ;
        RECT 94.430 -163.970 95.060 -160.120 ;
        RECT 96.450 -162.390 96.830 -161.710 ;
        RECT 117.190 -162.270 117.420 -161.810 ;
        RECT 96.985 -162.550 116.985 -162.320 ;
        RECT 97.160 -163.970 97.780 -162.550 ;
        RECT 88.040 -164.530 97.780 -163.970 ;
        RECT 88.040 -164.570 97.730 -164.530 ;
        RECT 88.040 -167.670 88.900 -164.570 ;
        RECT 94.430 -164.610 95.060 -164.570 ;
        RECT 68.970 -167.900 88.970 -167.670 ;
        RECT 68.460 -168.460 68.810 -167.920 ;
        RECT 89.130 -168.410 89.360 -167.950 ;
        RECT 66.290 -171.120 66.760 -171.080 ;
        RECT 63.660 -171.710 66.760 -171.120 ;
        RECT 68.820 -171.150 76.860 -171.140 ;
        RECT 68.730 -171.160 76.890 -171.150 ;
        RECT 68.730 -171.640 77.160 -171.160 ;
        RECT 63.660 -171.750 64.340 -171.710 ;
        RECT 66.290 -171.770 66.760 -171.710 ;
        RECT 74.500 -174.750 75.490 -174.650 ;
        RECT 74.100 -175.280 74.340 -174.890 ;
        RECT 74.490 -174.980 75.490 -174.750 ;
        RECT 75.630 -174.940 75.870 -174.850 ;
        RECT 75.630 -175.230 75.880 -174.940 ;
        RECT 75.630 -176.260 75.870 -175.230 ;
        RECT 76.880 -176.260 77.160 -171.640 ;
        RECT 78.880 -174.620 79.880 -174.610 ;
        RECT 78.840 -174.710 79.880 -174.620 ;
        RECT 78.400 -176.260 78.660 -174.830 ;
        RECT 78.835 -174.940 79.880 -174.710 ;
        RECT 80.070 -174.900 80.270 -174.840 ;
        RECT 78.840 -174.950 79.880 -174.940 ;
        RECT 80.040 -175.190 80.270 -174.900 ;
        RECT 80.070 -175.230 80.270 -175.190 ;
        RECT 75.630 -176.450 78.660 -176.260 ;
        RECT 75.610 -176.650 78.660 -176.450 ;
        RECT 75.610 -176.680 78.650 -176.650 ;
        RECT 75.610 -176.690 75.750 -176.680 ;
        RECT 76.880 -176.700 77.380 -176.680 ;
        RECT 62.640 -176.960 65.600 -176.950 ;
        RECT 77.130 -176.960 77.380 -176.700 ;
        RECT -2.320 -177.110 0.720 -177.080 ;
        RECT -2.320 -177.120 -2.180 -177.110 ;
        RECT -1.050 -177.130 -0.550 -177.110 ;
        RECT -15.290 -177.390 -12.330 -177.380 ;
        RECT -0.800 -177.390 -0.550 -177.130 ;
        RECT 62.640 -177.260 77.380 -176.960 ;
        RECT 62.640 -177.270 65.600 -177.260 ;
        RECT -15.290 -177.660 -0.550 -177.390 ;
        RECT 77.130 -177.320 77.380 -177.260 ;
        RECT 77.130 -177.440 77.440 -177.320 ;
        RECT -15.290 -177.690 -0.540 -177.660 ;
        RECT -15.290 -177.700 -12.330 -177.690 ;
        RECT -0.870 -182.740 -0.540 -177.690 ;
        RECT -0.910 -183.580 36.160 -182.740 ;
        RECT 35.500 -186.040 36.130 -183.580 ;
        RECT 33.690 -186.680 36.130 -186.040 ;
        RECT 33.690 -188.010 35.960 -186.680 ;
        RECT 33.430 -192.050 36.500 -188.010 ;
        RECT 47.300 -188.480 48.710 -188.420 ;
        RECT 77.150 -188.480 77.440 -177.440 ;
        RECT 47.300 -189.170 77.440 -188.480 ;
        RECT 47.300 -189.310 77.430 -189.170 ;
        RECT 47.300 -194.820 48.710 -189.310 ;
        RECT 46.250 -194.900 49.920 -194.820 ;
        RECT 46.210 -195.050 49.920 -194.900 ;
        RECT 46.210 -196.550 46.540 -195.050 ;
        RECT 49.590 -196.490 49.920 -195.050 ;
        RECT 45.220 -197.050 45.500 -196.720 ;
        RECT 45.660 -196.780 46.660 -196.550 ;
        RECT 46.810 -197.140 47.190 -196.580 ;
        RECT 49.030 -197.090 49.370 -196.590 ;
        RECT 49.565 -196.720 50.565 -196.490 ;
        RECT 50.760 -196.990 51.040 -196.660 ;
        RECT 47.940 -200.300 48.210 -200.290 ;
        RECT 47.940 -200.600 49.900 -200.300 ;
        RECT 45.680 -202.130 46.680 -201.900 ;
        RECT 46.230 -204.920 46.520 -202.130 ;
        RECT 47.940 -202.290 48.210 -200.600 ;
        RECT 49.680 -201.480 49.900 -200.600 ;
        RECT 49.495 -201.710 50.495 -201.480 ;
        RECT 47.900 -203.040 48.210 -202.290 ;
        RECT 47.900 -203.980 48.720 -203.040 ;
        RECT 45.790 -205.150 46.790 -204.920 ;
        RECT 45.790 -205.590 46.790 -205.360 ;
        RECT 46.400 -206.500 46.660 -205.590 ;
        RECT 47.900 -205.660 48.210 -203.980 ;
        RECT 49.475 -205.570 50.475 -205.340 ;
        RECT 47.900 -206.500 48.170 -205.660 ;
        RECT 46.400 -206.860 48.170 -206.500 ;
        RECT 46.400 -206.870 46.660 -206.860 ;
        RECT 47.900 -207.350 48.170 -206.860 ;
        RECT 49.620 -207.350 49.760 -205.570 ;
        RECT 47.900 -207.590 49.760 -207.350 ;
        RECT 47.900 -207.620 49.740 -207.590 ;
        RECT 47.900 -207.660 48.170 -207.620 ;
        RECT 47.670 -215.110 48.910 -213.700 ;
        RECT 46.090 -215.190 49.760 -215.110 ;
        RECT 46.050 -215.340 49.760 -215.190 ;
        RECT 46.050 -216.840 46.380 -215.340 ;
        RECT 49.430 -216.780 49.760 -215.340 ;
        RECT 45.060 -217.340 45.340 -217.010 ;
        RECT 45.500 -217.070 46.500 -216.840 ;
        RECT 46.650 -217.430 47.030 -216.870 ;
        RECT 48.870 -217.380 49.210 -216.880 ;
        RECT 49.405 -217.010 50.405 -216.780 ;
        RECT 50.600 -217.280 50.880 -216.950 ;
        RECT 47.780 -220.590 48.050 -220.580 ;
        RECT 47.780 -220.890 49.740 -220.590 ;
        RECT 45.520 -222.420 46.520 -222.190 ;
        RECT 46.070 -225.210 46.360 -222.420 ;
        RECT 47.780 -222.580 48.050 -220.890 ;
        RECT 49.520 -221.770 49.740 -220.890 ;
        RECT 49.335 -222.000 50.335 -221.770 ;
        RECT 47.740 -223.330 48.050 -222.580 ;
        RECT 47.740 -224.270 48.560 -223.330 ;
        RECT 45.170 -225.400 45.460 -225.380 ;
        RECT 45.170 -225.690 45.470 -225.400 ;
        RECT 45.630 -225.440 46.630 -225.210 ;
        RECT 45.170 -225.710 45.460 -225.690 ;
        RECT 45.210 -227.920 45.460 -225.710 ;
        RECT 45.630 -225.880 46.630 -225.650 ;
        RECT 46.780 -225.710 47.060 -225.380 ;
        RECT 46.240 -226.790 46.500 -225.880 ;
        RECT 47.740 -225.950 48.050 -224.270 ;
        RECT 50.530 -225.350 50.840 -225.340 ;
        RECT 48.820 -225.380 49.100 -225.350 ;
        RECT 48.820 -225.670 49.110 -225.380 ;
        RECT 48.820 -225.680 49.100 -225.670 ;
        RECT 49.315 -225.860 50.315 -225.630 ;
        RECT 50.500 -225.680 50.840 -225.350 ;
        RECT 47.740 -226.790 48.010 -225.950 ;
        RECT 46.240 -227.150 48.010 -226.790 ;
        RECT 46.240 -227.160 46.500 -227.150 ;
        RECT 45.200 -228.420 45.460 -227.920 ;
        RECT 47.740 -227.640 48.010 -227.150 ;
        RECT 49.460 -227.640 49.600 -225.860 ;
        RECT 47.740 -227.880 49.600 -227.640 ;
        RECT 47.740 -227.910 49.580 -227.880 ;
        RECT 47.740 -227.950 48.010 -227.910 ;
        RECT 45.200 -229.080 45.450 -228.420 ;
        RECT 50.530 -229.080 50.840 -225.680 ;
        RECT 45.200 -229.630 50.850 -229.080 ;
        RECT 47.590 -230.430 48.140 -229.630 ;
        RECT 46.920 -230.870 48.160 -230.430 ;
        RECT 46.920 -234.980 47.200 -230.870 ;
        RECT 45.230 -235.210 48.500 -234.980 ;
        RECT 45.230 -236.600 45.500 -235.210 ;
        RECT 48.240 -236.550 48.500 -235.210 ;
        RECT 44.600 -236.830 45.600 -236.600 ;
        RECT 47.965 -236.780 48.965 -236.550 ;
      LAYER via ;
        RECT 45.740 197.610 46.020 198.270 ;
        RECT 44.280 191.160 44.540 191.470 ;
        RECT 46.530 191.100 46.790 191.400 ;
        RECT 45.660 188.390 45.980 189.000 ;
        RECT 45.900 177.320 46.180 177.980 ;
        RECT 44.440 170.870 44.700 171.180 ;
        RECT 46.690 170.810 46.950 171.110 ;
        RECT 32.370 163.500 33.120 164.800 ;
        RECT -5.820 149.230 -4.860 149.490 ;
        RECT -1.460 149.210 -0.500 149.490 ;
        RECT -13.960 145.790 -13.700 146.100 ;
        RECT -11.450 145.790 -11.190 146.090 ;
        RECT -11.830 142.510 -11.570 142.980 ;
        RECT -13.960 138.650 -13.700 139.190 ;
        RECT -11.860 138.690 -11.590 139.100 ;
        RECT 16.160 136.330 16.420 136.860 ;
        RECT 14.240 132.560 14.850 133.080 ;
        RECT -11.830 130.310 -11.570 130.770 ;
        RECT 72.110 148.800 73.070 149.060 ;
        RECT 76.470 148.780 77.430 149.060 ;
        RECT 63.970 145.360 64.230 145.670 ;
        RECT 66.480 145.360 66.740 145.660 ;
        RECT 66.100 142.080 66.360 142.550 ;
        RECT 63.970 138.220 64.230 138.760 ;
        RECT 66.070 138.260 66.340 138.670 ;
        RECT 94.090 135.900 94.350 136.430 ;
        RECT 92.170 132.130 92.780 132.650 ;
        RECT 66.100 129.880 66.360 130.340 ;
        RECT 15.640 121.480 16.330 121.900 ;
        RECT 93.570 121.050 94.260 121.470 ;
        RECT 14.120 115.560 14.480 116.190 ;
        RECT 18.480 115.240 18.870 116.040 ;
        RECT 18.560 105.180 18.920 105.660 ;
        RECT 63.660 87.340 63.920 87.640 ;
        RECT -2.840 82.430 -2.580 82.700 ;
        RECT 63.890 83.690 64.150 83.950 ;
        RECT 62.540 82.120 62.800 82.460 ;
        RECT -222.270 40.540 -221.960 40.800 ;
        RECT -215.360 40.540 -214.820 40.800 ;
        RECT -219.150 38.410 -218.680 38.670 ;
        RECT -215.270 38.430 -214.860 38.700 ;
        RECT -206.940 38.410 -206.480 38.670 ;
        RECT -9.520 39.050 -8.970 39.760 ;
        RECT -222.260 38.030 -221.960 38.290 ;
        RECT -225.660 31.700 -225.400 32.660 ;
        RECT -240.970 -6.280 -239.670 -5.530 ;
        RECT -225.660 27.340 -225.380 28.300 ;
        RECT -115.930 35.810 -115.220 36.360 ;
        RECT 13.620 61.220 14.360 62.040 ;
        RECT 65.520 40.390 65.780 40.650 ;
        RECT -3.840 31.880 -3.560 32.250 ;
        RECT 0.730 33.620 0.990 33.880 ;
        RECT 65.560 36.590 65.820 36.850 ;
        RECT 64.140 34.740 64.530 35.360 ;
        RECT -108.420 30.400 -108.050 30.680 ;
        RECT -209.250 11.990 -208.730 12.600 ;
        RECT -158.870 29.420 -158.600 29.680 ;
        RECT 63.930 28.500 64.340 29.100 ;
        RECT -192.360 12.360 -191.730 12.720 ;
        RECT -213.030 10.420 -212.500 10.680 ;
        RECT -198.070 10.510 -197.650 11.200 ;
        RECT -192.210 7.970 -191.410 8.360 ;
        RECT -181.830 7.920 -181.350 8.280 ;
        RECT -138.210 12.480 -137.390 13.220 ;
        RECT -110.050 25.850 -109.790 26.110 ;
        RECT -1.320 3.820 -1.060 4.080 ;
        RECT -1.400 0.500 -1.140 0.760 ;
        RECT -267.640 -17.700 -267.330 -17.440 ;
        RECT -274.440 -19.180 -273.780 -18.900 ;
        RECT -247.350 -17.860 -247.040 -17.600 ;
        RECT -265.170 -19.140 -264.560 -18.820 ;
        RECT -267.570 -19.950 -267.270 -19.690 ;
        RECT -254.150 -19.340 -253.490 -19.060 ;
        RECT -247.280 -20.110 -246.980 -19.850 ;
        RECT -221.840 -37.390 -221.530 -37.130 ;
        RECT -214.930 -37.390 -214.390 -37.130 ;
        RECT -218.720 -39.520 -218.250 -39.260 ;
        RECT -214.840 -39.500 -214.430 -39.230 ;
        RECT -158.630 -35.960 -158.290 -35.700 ;
        RECT -163.810 -37.080 -163.510 -36.820 ;
        RECT -206.510 -39.520 -206.050 -39.260 ;
        RECT -160.120 -37.310 -159.860 -37.050 ;
        RECT -111.530 -37.690 -110.910 -37.300 ;
        RECT -105.270 -37.500 -104.670 -37.090 ;
        RECT -221.830 -39.900 -221.530 -39.640 ;
        RECT -225.230 -46.230 -224.970 -45.270 ;
        RECT -225.230 -50.590 -224.950 -49.630 ;
        RECT -116.820 -38.940 -116.560 -38.680 ;
        RECT -208.820 -65.940 -208.300 -65.330 ;
        RECT -113.020 -38.980 -112.760 -38.720 ;
        RECT -1.700 -45.240 -1.210 -44.930 ;
        RECT 66.450 -45.700 66.710 -45.440 ;
        RECT 66.350 -54.990 66.760 -54.390 ;
        RECT -1.420 -58.140 -1.140 -57.770 ;
        RECT -7.100 -65.650 -6.550 -64.940 ;
        RECT -212.600 -67.510 -212.070 -67.250 ;
        RECT -197.640 -67.420 -197.220 -66.730 ;
        RECT 3.150 -59.770 3.410 -59.510 ;
        RECT 66.560 -61.250 66.950 -60.630 ;
        RECT 67.980 -62.740 68.240 -62.480 ;
        RECT 67.940 -66.540 68.200 -66.280 ;
        RECT 16.040 -87.930 16.780 -87.110 ;
        RECT -0.420 -108.590 -0.160 -108.320 ;
        RECT 64.960 -108.350 65.220 -108.010 ;
        RECT 66.310 -109.840 66.570 -109.580 ;
        RECT 66.080 -113.530 66.340 -113.230 ;
        RECT 20.980 -131.550 21.340 -131.070 ;
        RECT 16.540 -142.080 16.900 -141.450 ;
        RECT 20.900 -141.930 21.290 -141.130 ;
        RECT 18.060 -147.790 18.750 -147.370 ;
        RECT 95.990 -147.360 96.680 -146.940 ;
        RECT -9.410 -156.660 -9.150 -156.200 ;
        RECT 16.660 -158.970 17.270 -158.450 ;
        RECT -11.540 -165.080 -11.280 -164.540 ;
        RECT -9.440 -164.990 -9.170 -164.580 ;
        RECT 18.580 -162.750 18.840 -162.220 ;
        RECT -9.410 -168.870 -9.150 -168.400 ;
        RECT -11.540 -171.990 -11.280 -171.680 ;
        RECT -9.030 -171.980 -8.770 -171.680 ;
        RECT -3.400 -175.380 -2.440 -175.120 ;
        RECT 0.960 -175.380 1.920 -175.100 ;
        RECT 68.520 -156.230 68.780 -155.770 ;
        RECT 94.590 -158.540 95.200 -158.020 ;
        RECT 66.390 -164.650 66.650 -164.110 ;
        RECT 68.490 -164.560 68.760 -164.150 ;
        RECT 96.510 -162.320 96.770 -161.790 ;
        RECT 68.520 -168.440 68.780 -167.970 ;
        RECT 66.390 -171.560 66.650 -171.250 ;
        RECT 68.900 -171.550 69.160 -171.250 ;
        RECT 74.530 -174.950 75.490 -174.690 ;
        RECT 78.890 -174.950 79.850 -174.670 ;
        RECT 34.790 -190.690 35.540 -189.390 ;
        RECT 46.860 -197.070 47.120 -196.760 ;
        RECT 49.110 -197.000 49.370 -196.700 ;
        RECT 48.320 -203.870 48.600 -203.210 ;
        RECT 48.080 -214.890 48.400 -214.280 ;
        RECT 46.700 -217.360 46.960 -217.050 ;
        RECT 48.950 -217.290 49.210 -216.990 ;
        RECT 48.160 -224.160 48.440 -223.500 ;
      LAYER met2 ;
        RECT 45.670 198.330 46.090 198.350 ;
        RECT 46.450 198.330 46.650 198.360 ;
        RECT 45.670 197.520 46.650 198.330 ;
        RECT 45.670 197.480 46.090 197.520 ;
        RECT 46.450 192.770 46.650 197.520 ;
        RECT 45.220 192.420 46.660 192.770 ;
        RECT 44.230 191.490 44.550 191.500 ;
        RECT 45.200 191.490 45.490 192.420 ;
        RECT 44.230 191.450 45.490 191.490 ;
        RECT 44.230 191.140 46.800 191.450 ;
        RECT 44.230 191.070 44.550 191.140 ;
        RECT 45.200 190.970 46.800 191.140 ;
        RECT 45.200 190.950 45.490 190.970 ;
        RECT 32.120 189.300 46.140 189.310 ;
        RECT 32.000 189.250 46.140 189.300 ;
        RECT 32.000 188.270 46.440 189.250 ;
        RECT 32.000 188.160 32.860 188.270 ;
        RECT 32.000 166.000 32.740 188.160 ;
        RECT 45.830 178.040 46.250 178.060 ;
        RECT 46.610 178.040 46.810 178.070 ;
        RECT 45.830 177.230 46.810 178.040 ;
        RECT 45.830 177.190 46.250 177.230 ;
        RECT 46.610 172.480 46.810 177.230 ;
        RECT 45.380 172.130 46.820 172.480 ;
        RECT 44.390 171.200 44.710 171.210 ;
        RECT 45.360 171.200 45.650 172.130 ;
        RECT 44.390 171.160 45.650 171.200 ;
        RECT 44.390 170.850 46.960 171.160 ;
        RECT 44.390 170.780 44.710 170.850 ;
        RECT 45.360 170.680 46.960 170.850 ;
        RECT 45.360 170.660 45.650 170.680 ;
        RECT 32.000 165.550 32.760 166.000 ;
        RECT 33.390 165.550 33.660 165.690 ;
        RECT 32.000 164.160 33.660 165.550 ;
        RECT 32.020 162.590 33.660 164.160 ;
        RECT -3.180 149.490 -2.960 149.510 ;
        RECT -5.960 149.230 -0.470 149.490 ;
        RECT -4.890 149.210 -0.470 149.230 ;
        RECT -14.840 147.600 -14.330 147.610 ;
        RECT -3.180 147.600 -2.960 149.210 ;
        RECT 74.750 149.060 74.970 149.080 ;
        RECT 71.970 148.800 77.460 149.060 ;
        RECT 73.040 148.780 77.460 148.800 ;
        RECT -14.840 147.190 -2.960 147.600 ;
        RECT -14.840 143.080 -14.330 147.190 ;
        RECT 63.090 147.170 63.600 147.180 ;
        RECT 74.750 147.170 74.970 148.780 ;
        RECT 63.090 146.760 74.970 147.170 ;
        RECT -11.670 146.190 -11.150 146.410 ;
        RECT -14.070 145.700 -11.150 146.190 ;
        RECT -13.860 145.690 -11.150 145.700 ;
        RECT -11.670 145.570 -11.150 145.690 ;
        RECT -11.940 143.080 -11.510 143.090 ;
        RECT -14.840 142.440 -11.510 143.080 ;
        RECT -14.840 133.670 -14.330 142.440 ;
        RECT -11.940 142.390 -11.510 142.440 ;
        RECT 63.090 142.650 63.600 146.760 ;
        RECT 66.260 145.760 66.780 145.980 ;
        RECT 63.860 145.270 66.780 145.760 ;
        RECT 64.070 145.260 66.780 145.270 ;
        RECT 66.260 145.140 66.780 145.260 ;
        RECT 65.990 142.650 66.420 142.660 ;
        RECT 63.090 142.010 66.420 142.650 ;
        RECT -14.040 139.240 -13.680 139.300 ;
        RECT -14.040 138.550 -11.560 139.240 ;
        RECT -14.040 138.490 -13.680 138.550 ;
        RECT -14.840 133.180 -11.490 133.670 ;
        RECT 13.970 133.200 14.990 133.280 ;
        RECT -14.330 133.170 -11.490 133.180 ;
        RECT -11.830 130.800 -11.590 133.170 ;
        RECT 13.780 132.310 14.990 133.200 ;
        RECT -11.860 130.280 -11.570 130.800 ;
        RECT 13.780 116.820 14.940 132.310 ;
        RECT 15.400 121.180 16.440 136.910 ;
        RECT 63.090 133.240 63.600 142.010 ;
        RECT 65.990 141.960 66.420 142.010 ;
        RECT 63.890 138.810 64.250 138.870 ;
        RECT 63.890 138.120 66.370 138.810 ;
        RECT 63.890 138.060 64.250 138.120 ;
        RECT 63.090 132.750 66.440 133.240 ;
        RECT 91.900 132.770 92.920 132.850 ;
        RECT 63.600 132.740 66.440 132.750 ;
        RECT 66.100 130.370 66.340 132.740 ;
        RECT 91.710 131.880 92.920 132.770 ;
        RECT 66.070 129.850 66.360 130.370 ;
        RECT 13.720 115.740 14.940 116.820 ;
        RECT 15.640 116.610 16.390 121.180 ;
        RECT 15.640 116.130 19.410 116.610 ;
        RECT 15.860 116.120 19.410 116.130 ;
        RECT 13.720 114.830 14.820 115.740 ;
        RECT 18.100 114.170 19.290 116.120 ;
        RECT 91.710 115.310 92.870 131.880 ;
        RECT 93.330 120.750 94.370 136.480 ;
        RECT 93.570 116.040 94.320 120.750 ;
        RECT 93.570 115.700 94.520 116.040 ;
        RECT 18.060 104.520 19.510 106.080 ;
        RECT -6.220 103.390 -5.570 103.450 ;
        RECT 18.450 103.390 18.970 104.520 ;
        RECT 91.820 104.240 92.700 115.310 ;
        RECT 61.170 104.180 92.800 104.240 ;
        RECT -6.220 102.570 19.030 103.390 ;
        RECT 61.030 103.030 92.800 104.180 ;
        RECT -6.220 82.980 -5.570 102.570 ;
        RECT -6.240 82.920 -5.570 82.980 ;
        RECT 52.730 87.690 53.330 87.800 ;
        RECT 61.030 87.720 61.610 103.030 ;
        RECT 63.540 87.720 63.950 87.940 ;
        RECT 61.030 87.690 63.950 87.720 ;
        RECT 52.730 87.290 63.950 87.690 ;
        RECT -6.250 82.140 -2.550 82.920 ;
        RECT -6.240 77.690 -5.950 82.140 ;
        RECT 13.710 77.690 14.220 77.790 ;
        RECT -6.240 77.200 14.220 77.690 ;
        RECT -6.240 77.160 -5.950 77.200 ;
        RECT 13.710 63.060 14.220 77.200 ;
        RECT 12.820 59.930 15.420 63.060 ;
        RECT -223.780 41.170 -209.350 41.680 ;
        RECT -225.660 31.730 -225.400 32.800 ;
        RECT -225.660 30.020 -225.380 31.730 ;
        RECT -223.770 30.020 -223.360 41.170 ;
        RECT -222.360 40.700 -221.870 40.910 ;
        RECT -222.360 38.510 -221.860 40.700 ;
        RECT -219.250 38.780 -218.610 41.170 ;
        RECT -215.470 40.520 -214.660 40.880 ;
        RECT -222.580 37.990 -221.740 38.510 ;
        RECT -219.260 38.350 -218.560 38.780 ;
        RECT -215.410 38.400 -214.720 40.520 ;
        RECT -209.840 38.670 -209.340 41.170 ;
        RECT -10.030 39.830 -8.340 40.280 ;
        RECT -10.030 39.160 -0.400 39.830 ;
        RECT -206.970 38.670 -206.450 38.700 ;
        RECT -209.840 38.430 -206.450 38.670 ;
        RECT -209.840 38.330 -209.340 38.430 ;
        RECT -206.970 38.410 -206.450 38.430 ;
        RECT -10.030 38.180 -8.340 39.160 ;
        RECT -116.450 35.180 -114.350 36.870 ;
        RECT -159.090 33.080 -158.310 33.090 ;
        RECT -159.150 33.060 -153.330 33.080 ;
        RECT -179.620 32.790 -153.330 33.060 ;
        RECT -179.620 32.410 -158.310 32.790 ;
        RECT -225.680 29.800 -223.360 30.020 ;
        RECT -225.660 27.310 -225.380 29.800 ;
        RECT -192.990 13.060 -191.000 13.120 ;
        RECT -209.370 12.870 -191.000 13.060 ;
        RECT -209.450 12.020 -191.000 12.870 ;
        RECT -209.450 11.900 -191.910 12.020 ;
        RECT -209.450 11.850 -208.480 11.900 ;
        RECT -213.080 11.200 -197.350 11.440 ;
        RECT -213.080 10.980 -192.300 11.200 ;
        RECT -213.080 10.450 -192.290 10.980 ;
        RECT -213.080 10.400 -197.350 10.450 ;
        RECT -192.780 8.740 -192.290 10.450 ;
        RECT -192.780 7.550 -190.340 8.740 ;
        RECT -182.250 8.390 -180.690 8.780 ;
        RECT -179.560 8.390 -178.740 32.410 ;
        RECT -159.090 29.390 -158.310 32.410 ;
        RECT -153.860 13.130 -153.370 32.790 ;
        RECT -116.000 27.420 -115.330 35.180 ;
        RECT -0.580 33.900 -0.400 39.160 ;
        RECT 0.620 33.900 1.020 34.120 ;
        RECT -0.580 33.600 1.020 33.900 ;
        RECT 0.620 33.260 1.020 33.600 ;
        RECT -4.250 31.280 -3.080 32.660 ;
        RECT -108.830 30.750 -107.450 31.090 ;
        RECT -95.740 30.750 -78.880 30.860 ;
        RECT -108.830 30.330 -78.880 30.750 ;
        RECT -108.830 29.920 -107.450 30.330 ;
        RECT -95.740 30.240 -78.880 30.330 ;
        RECT -116.000 27.240 -109.770 27.420 ;
        RECT -110.070 26.220 -109.770 27.240 ;
        RECT -110.290 25.820 -109.430 26.220 ;
        RECT -139.230 13.130 -136.100 14.020 ;
        RECT -153.960 12.620 -136.100 13.130 ;
        RECT -139.230 11.420 -136.100 12.620 ;
        RECT -182.250 7.870 -178.740 8.390 ;
        RECT -192.780 7.430 -192.290 7.550 ;
        RECT -182.250 7.330 -180.690 7.870 ;
        RECT -179.560 7.810 -178.740 7.870 ;
        RECT -79.590 3.870 -78.880 30.240 ;
        RECT -3.910 20.440 -3.490 31.280 ;
        RECT 52.730 30.010 53.330 87.290 ;
        RECT 61.030 87.270 63.950 87.290 ;
        RECT 61.030 87.080 61.610 87.270 ;
        RECT 63.540 86.950 63.950 87.270 ;
        RECT 63.630 83.500 64.250 84.230 ;
        RECT 62.370 81.890 63.000 82.620 ;
        RECT 62.460 38.830 62.880 81.890 ;
        RECT 63.740 73.460 64.240 83.500 ;
        RECT 63.740 73.370 64.910 73.460 ;
        RECT 93.590 73.370 94.520 115.700 ;
        RECT 63.740 72.450 94.520 73.370 ;
        RECT 63.740 72.260 94.230 72.450 ;
        RECT 63.740 72.220 64.910 72.260 ;
        RECT 63.920 72.180 64.910 72.220 ;
        RECT 65.400 40.930 65.680 72.260 ;
        RECT 65.380 40.000 65.810 40.930 ;
        RECT 62.460 37.900 62.970 38.830 ;
        RECT 62.460 37.730 62.920 37.900 ;
        RECT 62.510 35.360 62.920 37.730 ;
        RECT 65.410 36.250 65.870 37.120 ;
        RECT 63.740 35.360 65.020 35.880 ;
        RECT 62.510 34.690 65.020 35.360 ;
        RECT 62.510 34.580 62.920 34.690 ;
        RECT 63.740 33.790 65.020 34.690 ;
        RECT 54.750 31.010 55.320 31.050 ;
        RECT 65.540 31.010 65.860 36.250 ;
        RECT 54.750 30.610 65.890 31.010 ;
        RECT 54.750 30.010 55.320 30.610 ;
        RECT 52.730 29.450 55.320 30.010 ;
        RECT 52.750 29.340 55.320 29.450 ;
        RECT 54.750 29.300 55.320 29.340 ;
        RECT 63.410 27.610 64.980 29.600 ;
        RECT -3.970 19.220 -3.490 20.440 ;
        RECT 63.880 19.930 64.410 27.610 ;
        RECT -3.970 9.680 -3.540 19.220 ;
        RECT 3.310 9.680 3.960 9.690 ;
        RECT -4.010 9.090 4.060 9.680 ;
        RECT 3.310 7.990 3.960 9.090 ;
        RECT 63.770 8.280 64.500 19.930 ;
        RECT 3.350 6.440 3.940 7.990 ;
        RECT 7.420 7.870 64.860 8.280 ;
        RECT 7.450 7.200 8.040 7.870 ;
        RECT 7.430 7.090 8.040 7.200 ;
        RECT 7.430 6.475 8.020 7.090 ;
        RECT 3.335 5.030 3.940 6.440 ;
        RECT 3.335 4.770 3.470 5.030 ;
        RECT 3.730 4.770 3.940 5.030 ;
        RECT -1.520 3.890 -0.860 4.220 ;
        RECT -1.910 3.870 -0.860 3.890 ;
        RECT -79.590 3.630 -0.860 3.870 ;
        RECT 3.335 3.840 3.940 4.770 ;
        RECT 7.410 5.050 8.020 6.475 ;
        RECT 7.410 4.790 7.550 5.050 ;
        RECT 7.810 4.790 8.020 5.050 ;
        RECT 7.410 3.860 8.020 4.790 ;
        RECT -79.590 3.580 -1.060 3.630 ;
        RECT -79.590 3.470 -78.880 3.580 ;
        RECT -1.910 3.500 -1.060 3.580 ;
        RECT 3.335 3.000 3.905 3.840 ;
        RECT 7.410 3.020 7.980 3.860 ;
        RECT 3.300 1.590 3.905 3.000 ;
        RECT 3.300 1.330 3.430 1.590 ;
        RECT 3.690 1.330 3.905 1.590 ;
        RECT -1.610 0.290 -0.940 0.870 ;
        RECT 3.300 0.400 3.905 1.330 ;
        RECT 7.360 1.610 7.980 3.020 ;
        RECT 7.360 1.350 7.490 1.610 ;
        RECT 7.750 1.350 7.980 1.610 ;
        RECT 7.360 0.425 7.980 1.350 ;
        RECT 7.360 0.420 7.960 0.425 ;
        RECT 3.335 0.390 3.905 0.400 ;
        RECT -80.190 -3.070 -79.630 -2.900 ;
        RECT -80.430 -3.090 -3.030 -3.070 ;
        RECT -1.540 -3.090 -1.130 0.290 ;
        RECT -80.430 -3.360 -0.900 -3.090 ;
        RECT -265.470 -5.180 -240.330 -5.160 ;
        RECT -265.470 -5.280 -238.760 -5.180 ;
        RECT -265.480 -5.900 -238.760 -5.280 ;
        RECT -265.480 -6.020 -264.330 -5.900 ;
        RECT -242.170 -5.920 -238.760 -5.900 ;
        RECT -267.670 -17.710 -267.240 -17.390 ;
        RECT -267.660 -18.360 -267.310 -17.710 ;
        RECT -268.590 -18.380 -267.120 -18.360 ;
        RECT -268.940 -18.650 -267.120 -18.380 ;
        RECT -274.520 -19.250 -273.650 -18.830 ;
        RECT -274.500 -19.610 -273.690 -19.250 ;
        RECT -268.940 -19.610 -268.590 -18.650 ;
        RECT -274.530 -19.810 -268.590 -19.610 ;
        RECT -268.940 -19.820 -268.590 -19.810 ;
        RECT -267.620 -19.960 -267.140 -18.650 ;
        RECT -265.480 -19.300 -264.440 -6.020 ;
        RECT -241.720 -6.550 -238.760 -5.920 ;
        RECT -241.860 -6.820 -238.760 -6.550 ;
        RECT -247.380 -17.870 -246.950 -17.550 ;
        RECT -247.370 -18.520 -247.020 -17.870 ;
        RECT -248.300 -18.540 -246.830 -18.520 ;
        RECT -248.650 -18.810 -246.830 -18.540 ;
        RECT -265.420 -19.600 -264.440 -19.300 ;
        RECT -254.230 -19.410 -253.360 -18.990 ;
        RECT -254.210 -19.770 -253.400 -19.410 ;
        RECT -248.650 -19.770 -248.300 -18.810 ;
        RECT -254.240 -19.970 -248.300 -19.770 ;
        RECT -248.650 -19.980 -248.300 -19.970 ;
        RECT -247.330 -20.120 -246.850 -18.810 ;
        RECT -163.970 -25.910 -105.620 -25.890 ;
        RECT -163.970 -26.490 -105.510 -25.910 ;
        RECT -163.860 -34.190 -163.460 -26.490 ;
        RECT -106.180 -27.910 -105.510 -26.490 ;
        RECT -107.220 -28.480 -105.470 -27.910 ;
        RECT -180.350 -34.330 -163.250 -34.190 ;
        RECT -180.410 -34.770 -163.250 -34.330 ;
        RECT -223.350 -36.760 -208.920 -36.250 ;
        RECT -225.230 -46.200 -224.970 -45.130 ;
        RECT -225.230 -47.910 -224.950 -46.200 ;
        RECT -223.340 -47.910 -222.930 -36.760 ;
        RECT -221.930 -37.230 -221.440 -37.020 ;
        RECT -221.930 -39.420 -221.430 -37.230 ;
        RECT -218.820 -39.150 -218.180 -36.760 ;
        RECT -215.040 -37.410 -214.230 -37.050 ;
        RECT -222.150 -39.940 -221.310 -39.420 ;
        RECT -218.830 -39.580 -218.130 -39.150 ;
        RECT -214.980 -39.530 -214.290 -37.410 ;
        RECT -209.410 -39.260 -208.910 -36.760 ;
        RECT -206.540 -39.260 -206.020 -39.230 ;
        RECT -209.410 -39.500 -206.020 -39.260 ;
        RECT -209.410 -39.600 -208.910 -39.500 ;
        RECT -206.540 -39.520 -206.020 -39.500 ;
        RECT -225.250 -48.130 -222.930 -47.910 ;
        RECT -225.230 -50.620 -224.950 -48.130 ;
        RECT -208.940 -64.980 -191.480 -64.870 ;
        RECT -180.410 -64.980 -179.200 -34.770 ;
        RECT -163.890 -36.700 -163.440 -34.770 ;
        RECT -158.790 -35.620 -158.060 -35.530 ;
        RECT -158.790 -35.670 -113.900 -35.620 ;
        RECT -158.790 -36.040 -110.750 -35.670 ;
        RECT -158.790 -36.160 -158.060 -36.040 ;
        RECT -115.000 -36.080 -110.750 -36.040 ;
        RECT -115.000 -36.130 -114.070 -36.080 ;
        RECT -164.110 -37.110 -163.120 -36.700 ;
        RECT -160.400 -36.900 -159.670 -36.790 ;
        RECT -111.530 -36.900 -110.860 -36.080 ;
        RECT -160.400 -37.080 -148.390 -36.900 ;
        RECT -160.400 -37.400 -148.350 -37.080 ;
        RECT -160.400 -37.410 -159.670 -37.400 ;
        RECT -149.630 -38.070 -148.350 -37.400 ;
        RECT -208.940 -65.060 -179.200 -64.980 ;
        RECT -209.020 -65.860 -179.200 -65.060 ;
        RECT -209.020 -66.030 -191.480 -65.860 ;
        RECT -180.410 -65.960 -179.200 -65.860 ;
        RECT -149.540 -38.560 -148.430 -38.070 ;
        RECT -112.050 -38.180 -109.960 -36.900 ;
        RECT -117.100 -38.560 -116.170 -38.540 ;
        RECT -149.540 -38.840 -116.170 -38.560 ;
        RECT -209.020 -66.080 -208.050 -66.030 ;
        RECT -212.650 -66.730 -196.920 -66.490 ;
        RECT -212.650 -66.750 -191.870 -66.730 ;
        RECT -149.540 -66.750 -148.430 -38.840 ;
        RECT -117.100 -38.970 -116.170 -38.840 ;
        RECT -113.290 -38.700 -112.420 -38.570 ;
        RECT -107.180 -38.700 -106.780 -28.480 ;
        RECT -105.770 -37.040 -103.780 -36.570 ;
        RECT -105.770 -37.260 -95.760 -37.040 ;
        RECT -80.190 -37.250 -79.630 -3.360 ;
        RECT -3.180 -3.380 -0.900 -3.360 ;
        RECT -1.540 -3.410 -1.130 -3.380 ;
        RECT -90.680 -37.260 -79.630 -37.250 ;
        RECT -105.770 -37.570 -79.630 -37.260 ;
        RECT -105.770 -38.140 -103.780 -37.570 ;
        RECT -96.270 -37.620 -79.630 -37.570 ;
        RECT -90.680 -37.660 -79.630 -37.620 ;
        RECT -80.190 -37.900 -79.630 -37.660 ;
        RECT -113.290 -39.020 -106.780 -38.700 ;
        RECT -113.290 -39.030 -112.420 -39.020 ;
        RECT -107.180 -39.050 -106.780 -39.020 ;
        RECT -2.000 -45.480 -0.770 -44.570 ;
        RECT -1.490 -57.170 -1.070 -45.480 ;
        RECT 66.170 -45.890 67.030 -45.350 ;
        RECT 66.300 -53.500 66.830 -45.890 ;
        RECT 57.170 -55.230 57.740 -55.190 ;
        RECT 55.170 -55.340 57.740 -55.230 ;
        RECT 55.150 -55.900 57.740 -55.340 ;
        RECT 65.830 -55.490 67.400 -53.500 ;
        RECT -1.830 -58.550 -0.660 -57.170 ;
        RECT 3.040 -59.490 3.440 -59.150 ;
        RECT 1.840 -59.790 3.440 -59.490 ;
        RECT -7.610 -65.050 -5.920 -64.070 ;
        RECT 1.840 -65.050 2.020 -59.790 ;
        RECT 3.040 -60.010 3.440 -59.790 ;
        RECT -7.610 -65.720 2.020 -65.050 ;
        RECT -7.610 -66.170 -5.920 -65.720 ;
        RECT -212.650 -67.390 -148.430 -66.750 ;
        RECT -212.650 -67.480 -148.620 -67.390 ;
        RECT -212.650 -67.530 -196.920 -67.480 ;
        RECT -192.210 -67.680 -148.620 -67.480 ;
        RECT 15.240 -88.950 17.840 -85.820 ;
        RECT -3.820 -103.090 -3.530 -103.050 ;
        RECT 16.130 -103.090 16.640 -88.950 ;
        RECT -3.820 -103.580 16.640 -103.090 ;
        RECT -3.820 -108.030 -3.530 -103.580 ;
        RECT 16.130 -103.680 16.640 -103.580 ;
        RECT -3.830 -108.810 -0.130 -108.030 ;
        RECT -3.820 -108.870 -3.150 -108.810 ;
        RECT -3.800 -128.460 -3.150 -108.870 ;
        RECT 55.150 -113.180 55.750 -55.900 ;
        RECT 57.170 -56.500 57.740 -55.900 ;
        RECT 57.170 -56.900 68.310 -56.500 ;
        RECT 57.170 -56.940 57.740 -56.900 ;
        RECT 64.930 -60.580 65.340 -60.470 ;
        RECT 66.160 -60.580 67.440 -59.680 ;
        RECT 64.930 -61.250 67.440 -60.580 ;
        RECT 64.930 -63.620 65.340 -61.250 ;
        RECT 66.160 -61.770 67.440 -61.250 ;
        RECT 67.960 -62.140 68.280 -56.900 ;
        RECT 67.830 -63.010 68.290 -62.140 ;
        RECT 64.880 -63.790 65.340 -63.620 ;
        RECT 64.880 -64.720 65.390 -63.790 ;
        RECT 64.880 -107.780 65.300 -64.720 ;
        RECT 67.800 -66.820 68.230 -65.890 ;
        RECT 66.340 -98.110 67.330 -98.070 ;
        RECT 66.160 -98.150 67.330 -98.110 ;
        RECT 67.820 -98.150 68.100 -66.820 ;
        RECT 66.160 -98.340 96.650 -98.150 ;
        RECT 66.160 -99.260 96.940 -98.340 ;
        RECT 66.160 -99.350 67.330 -99.260 ;
        RECT 64.790 -108.510 65.420 -107.780 ;
        RECT 66.160 -109.390 66.660 -99.350 ;
        RECT 66.050 -110.120 66.670 -109.390 ;
        RECT 63.450 -113.160 64.030 -112.970 ;
        RECT 65.960 -113.160 66.370 -112.840 ;
        RECT 63.450 -113.180 66.370 -113.160 ;
        RECT 55.150 -113.580 66.370 -113.180 ;
        RECT 55.150 -113.690 55.750 -113.580 ;
        RECT 63.450 -113.610 66.370 -113.580 ;
        RECT -3.800 -129.280 21.450 -128.460 ;
        RECT 63.450 -128.920 64.030 -113.610 ;
        RECT 65.960 -113.830 66.370 -113.610 ;
        RECT -3.800 -129.340 -3.150 -129.280 ;
        RECT 20.870 -130.410 21.390 -129.280 ;
        RECT 63.450 -130.070 95.220 -128.920 ;
        RECT 63.590 -130.130 95.220 -130.070 ;
        RECT 20.480 -131.970 21.930 -130.410 ;
        RECT 16.140 -141.630 17.240 -140.720 ;
        RECT 16.140 -142.710 17.360 -141.630 ;
        RECT 20.520 -142.010 21.710 -140.060 ;
        RECT 94.240 -141.200 95.120 -130.130 ;
        RECT 18.280 -142.020 21.830 -142.010 ;
        RECT -9.440 -156.690 -9.150 -156.170 ;
        RECT -9.410 -159.060 -9.170 -156.690 ;
        RECT 16.200 -158.200 17.360 -142.710 ;
        RECT 18.060 -142.500 21.830 -142.020 ;
        RECT 18.060 -147.070 18.810 -142.500 ;
        RECT -11.910 -159.070 -9.070 -159.060 ;
        RECT -12.420 -159.560 -9.070 -159.070 ;
        RECT 16.200 -159.090 17.410 -158.200 ;
        RECT 16.390 -159.170 17.410 -159.090 ;
        RECT -12.420 -168.330 -11.910 -159.560 ;
        RECT 17.820 -162.800 18.860 -147.070 ;
        RECT 68.490 -156.260 68.780 -155.740 ;
        RECT 68.520 -158.630 68.760 -156.260 ;
        RECT 94.130 -157.770 95.290 -141.200 ;
        RECT 96.010 -141.590 96.940 -99.260 ;
        RECT 95.990 -141.930 96.940 -141.590 ;
        RECT 95.990 -146.640 96.740 -141.930 ;
        RECT 66.020 -158.640 68.860 -158.630 ;
        RECT 65.510 -159.130 68.860 -158.640 ;
        RECT 94.130 -158.660 95.340 -157.770 ;
        RECT 94.320 -158.740 95.340 -158.660 ;
        RECT -11.620 -164.440 -11.260 -164.380 ;
        RECT -11.620 -165.130 -9.140 -164.440 ;
        RECT -11.620 -165.190 -11.260 -165.130 ;
        RECT 65.510 -167.900 66.020 -159.130 ;
        RECT 95.750 -162.370 96.790 -146.640 ;
        RECT 66.310 -164.010 66.670 -163.950 ;
        RECT 66.310 -164.700 68.790 -164.010 ;
        RECT 66.310 -164.760 66.670 -164.700 ;
        RECT 68.410 -167.900 68.840 -167.850 ;
        RECT -9.520 -168.330 -9.090 -168.280 ;
        RECT -12.420 -168.970 -9.090 -168.330 ;
        RECT -12.420 -173.080 -11.910 -168.970 ;
        RECT -9.520 -168.980 -9.090 -168.970 ;
        RECT 65.510 -168.540 68.840 -167.900 ;
        RECT -9.250 -171.580 -8.730 -171.460 ;
        RECT -11.440 -171.590 -8.730 -171.580 ;
        RECT -11.650 -172.080 -8.730 -171.590 ;
        RECT -9.250 -172.300 -8.730 -172.080 ;
        RECT 65.510 -172.650 66.020 -168.540 ;
        RECT 68.410 -168.550 68.840 -168.540 ;
        RECT 68.680 -171.150 69.200 -171.030 ;
        RECT 66.490 -171.160 69.200 -171.150 ;
        RECT 66.280 -171.650 69.200 -171.160 ;
        RECT 68.680 -171.870 69.200 -171.650 ;
        RECT 65.510 -173.060 77.390 -172.650 ;
        RECT 65.510 -173.070 66.020 -173.060 ;
        RECT -12.420 -173.490 -0.540 -173.080 ;
        RECT -12.420 -173.500 -11.910 -173.490 ;
        RECT -0.760 -175.100 -0.540 -173.490 ;
        RECT 77.170 -174.670 77.390 -173.060 ;
        RECT 75.460 -174.690 79.880 -174.670 ;
        RECT 74.390 -174.950 79.880 -174.690 ;
        RECT 77.170 -174.970 77.390 -174.950 ;
        RECT -2.470 -175.120 1.950 -175.100 ;
        RECT -3.540 -175.380 1.950 -175.120 ;
        RECT -0.760 -175.400 -0.540 -175.380 ;
        RECT 34.440 -190.050 36.080 -188.480 ;
        RECT 34.420 -191.440 36.080 -190.050 ;
        RECT 34.420 -191.890 35.180 -191.440 ;
        RECT 35.810 -191.580 36.080 -191.440 ;
        RECT 34.420 -214.050 35.160 -191.890 ;
        RECT 47.780 -196.570 48.070 -196.550 ;
        RECT 46.810 -196.740 47.130 -196.670 ;
        RECT 47.780 -196.740 49.380 -196.570 ;
        RECT 46.810 -197.050 49.380 -196.740 ;
        RECT 46.810 -197.090 48.070 -197.050 ;
        RECT 46.810 -197.100 47.130 -197.090 ;
        RECT 47.780 -198.020 48.070 -197.090 ;
        RECT 47.800 -198.370 49.240 -198.020 ;
        RECT 48.250 -203.120 48.670 -203.080 ;
        RECT 49.030 -203.120 49.230 -198.370 ;
        RECT 48.250 -203.930 49.230 -203.120 ;
        RECT 48.250 -203.950 48.670 -203.930 ;
        RECT 49.030 -203.960 49.230 -203.930 ;
        RECT 34.420 -214.160 35.280 -214.050 ;
        RECT 34.420 -215.140 48.860 -214.160 ;
        RECT 34.420 -215.190 48.560 -215.140 ;
        RECT 34.540 -215.200 48.560 -215.190 ;
        RECT 47.620 -216.860 47.910 -216.840 ;
        RECT 46.650 -217.030 46.970 -216.960 ;
        RECT 47.620 -217.030 49.220 -216.860 ;
        RECT 46.650 -217.340 49.220 -217.030 ;
        RECT 46.650 -217.380 47.910 -217.340 ;
        RECT 46.650 -217.390 46.970 -217.380 ;
        RECT 47.620 -218.310 47.910 -217.380 ;
        RECT 47.640 -218.660 49.080 -218.310 ;
        RECT 48.090 -223.410 48.510 -223.370 ;
        RECT 48.870 -223.410 49.070 -218.660 ;
        RECT 48.090 -224.220 49.070 -223.410 ;
        RECT 48.090 -224.240 48.510 -224.220 ;
        RECT 48.870 -224.250 49.070 -224.220 ;
  END
END core_flat_v4
END LIBRARY

