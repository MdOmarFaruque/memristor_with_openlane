VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO core_flat_v4
  CLASS BLOCK ;
  FOREIGN core_flat_v4 ;
  ORIGIN 400.160 350.900 ;
  SIZE 650.010 BY 679.000 ;
  PIN SEL1
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT -400.160 -17.780 -398.160 -17.180 ;
    END
  END SEL1
  PIN DIGITALIN1
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT -400.130 -19.850 -398.160 -19.250 ;
    END
  END DIGITALIN1
  PIN AIN1
    ANTENNADIFFAREA 23.199999 ;
    PORT
      LAYER met3 ;
        RECT -400.160 -13.070 -398.160 -12.470 ;
    END
  END AIN1
  PIN SEL3
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 46.690 -350.900 46.990 -348.900 ;
    END
  END SEL3
  PIN DIGITALIN3
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 50.250 -350.890 50.550 -348.900 ;
    END
  END DIGITALIN3
  PIN AIN3
    ANTENNADIFFAREA 23.199999 ;
    PORT
      LAYER met2 ;
        RECT 41.840 -350.900 42.140 -348.900 ;
    END
  END AIN3
  PIN SEL2
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 44.330 326.100 44.630 328.100 ;
    END
  END SEL2
  PIN DIGITALIN2
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 47.090 326.100 47.390 328.090 ;
    END
  END DIGITALIN2
  PIN AIN2
    ANTENNADIFFAREA 23.199999 ;
    PORT
      LAYER met2 ;
        RECT 39.740 326.100 40.040 328.100 ;
    END
  END AIN2
  PIN vssa1
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT -400.150 241.100 249.850 251.100 ;
        RECT -400.150 -273.900 -398.160 -263.900 ;
        RECT 247.850 -273.900 249.850 -263.900 ;
    END
  END vssa1
  PIN vdda1
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT -400.150 266.100 -398.160 276.100 ;
        RECT 247.850 266.100 249.850 276.100 ;
        RECT -400.150 -298.900 249.850 -288.900 ;
    END
  END vdda1
  PIN vssd1
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT -400.150 291.100 -398.160 301.100 ;
        RECT 247.850 291.100 249.850 301.100 ;
        RECT -400.150 -323.900 249.850 -313.900 ;
    END
  END vssd1
  PIN vccd1
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT -252.750 -348.940 -252.270 -348.900 ;
      LAYER met3 ;
        RECT -400.150 316.100 -398.160 326.100 ;
        RECT 247.850 316.100 249.850 326.100 ;
        RECT -400.150 -348.900 249.850 -338.900 ;
    END
  END vccd1
  OBS
      LAYER li1 ;
        RECT -288.090 -237.810 118.140 211.920 ;
      LAYER met1 ;
        RECT -299.830 -256.200 151.420 233.660 ;
      LAYER met2 ;
        RECT -390.150 -348.900 239.850 326.100 ;
      LAYER met3 ;
        RECT -398.160 -273.900 247.850 326.100 ;
  END
END core_flat_v4
END LIBRARY

