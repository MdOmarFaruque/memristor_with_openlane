magic
tech sky130B
magscale 1 2
timestamp 1713777132
<< checkpaint >>
rect -12658 -11586 596582 715522
<< metal1 >>
rect 115106 1300 115112 1352
rect 115164 1340 115170 1352
rect 579614 1340 579620 1352
rect 115164 1312 579620 1340
rect 115164 1300 115170 1312
rect 579614 1300 579620 1312
rect 579672 1300 579678 1352
rect 244274 1232 244280 1284
rect 244332 1272 244338 1284
rect 580350 1272 580356 1284
rect 244332 1244 580356 1272
rect 244332 1232 244338 1244
rect 580350 1232 580356 1244
rect 580408 1232 580414 1284
rect 262858 1164 262864 1216
rect 262916 1204 262922 1216
rect 580534 1204 580540 1216
rect 262916 1176 580540 1204
rect 262916 1164 262922 1176
rect 580534 1164 580540 1176
rect 580592 1164 580598 1216
rect 282178 1096 282184 1148
rect 282236 1136 282242 1148
rect 580626 1136 580632 1148
rect 282236 1108 580632 1136
rect 282236 1096 282242 1108
rect 580626 1096 580632 1108
rect 580684 1096 580690 1148
rect 224954 620 224960 672
rect 225012 660 225018 672
rect 580350 660 580356 672
rect 225012 632 580356 660
rect 225012 620 225018 632
rect 580350 620 580356 632
rect 580408 620 580414 672
<< via1 >>
rect 115112 1300 115164 1352
rect 579620 1300 579672 1352
rect 244280 1232 244332 1284
rect 580356 1232 580408 1284
rect 262864 1164 262916 1216
rect 580540 1164 580592 1216
rect 282184 1096 282236 1148
rect 580632 1096 580684 1148
rect 224960 620 225012 672
rect 580356 620 580408 672
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 1193 8156 703520
rect 56796 700641 56824 703520
rect 12070 700632 12126 700641
rect 12070 700567 12126 700576
rect 56782 700632 56838 700641
rect 56782 700567 56838 700576
rect 9586 700360 9642 700369
rect 9586 700295 9642 700304
rect 9600 236201 9628 700295
rect 9586 236192 9642 236201
rect 9586 236127 9642 236136
rect 12084 49881 12112 700567
rect 12254 700496 12310 700505
rect 12254 700431 12310 700440
rect 12162 281480 12218 281489
rect 12162 281415 12218 281424
rect 12070 49872 12126 49881
rect 12070 49807 12126 49816
rect 12176 3369 12204 281415
rect 12268 143449 12296 700431
rect 71778 531312 71834 531321
rect 71778 531247 71834 531256
rect 71792 524498 71820 531247
rect 71700 524470 71820 524498
rect 71700 523025 71728 524470
rect 66902 523016 66958 523025
rect 66902 522951 66958 522960
rect 71686 523016 71742 523025
rect 71686 522951 71742 522960
rect 66916 506569 66944 522951
rect 65522 506560 65578 506569
rect 65522 506495 65578 506504
rect 66902 506560 66958 506569
rect 66902 506495 66958 506504
rect 65536 487393 65564 506495
rect 65522 487384 65578 487393
rect 65522 487319 65578 487328
rect 62762 487112 62818 487121
rect 62762 487047 62818 487056
rect 62776 475425 62804 487047
rect 60738 475416 60794 475425
rect 60738 475351 60794 475360
rect 62762 475416 62818 475425
rect 62762 475351 62818 475360
rect 60752 473362 60780 475351
rect 60660 473334 60780 473362
rect 60660 473249 60688 473334
rect 58622 473240 58678 473249
rect 58622 473175 58678 473184
rect 60646 473240 60702 473249
rect 60646 473175 60702 473184
rect 58636 459649 58664 473175
rect 56874 459640 56930 459649
rect 56874 459575 56930 459584
rect 58622 459640 58678 459649
rect 58622 459575 58678 459584
rect 56888 458289 56916 459575
rect 54482 458280 54538 458289
rect 54482 458215 54538 458224
rect 56874 458280 56930 458289
rect 56874 458215 56930 458224
rect 54496 446457 54524 458215
rect 53102 446448 53158 446457
rect 53102 446383 53158 446392
rect 54482 446448 54538 446457
rect 54482 446383 54538 446392
rect 53116 434761 53144 446383
rect 53102 434752 53158 434761
rect 53102 434687 53158 434696
rect 46938 434616 46994 434625
rect 46938 434551 46994 434560
rect 46952 427938 46980 434551
rect 46860 427910 46980 427938
rect 46860 422385 46888 427910
rect 42798 422376 42854 422385
rect 42798 422311 42854 422320
rect 46846 422376 46902 422385
rect 46846 422311 46902 422320
rect 42812 421002 42840 422311
rect 42720 420974 42840 421002
rect 42720 418305 42748 420974
rect 38566 418296 38622 418305
rect 38566 418231 38622 418240
rect 42706 418296 42762 418305
rect 42706 418231 42762 418240
rect 38580 412729 38608 418231
rect 38566 412720 38622 412729
rect 38566 412655 38622 412664
rect 31758 412584 31814 412593
rect 31758 412519 31814 412528
rect 31772 408921 31800 412519
rect 72988 409193 73016 703520
rect 121656 700505 121684 703520
rect 121642 700496 121698 700505
rect 121642 700431 121698 700440
rect 137848 699825 137876 703520
rect 186516 700369 186544 703520
rect 186502 700360 186558 700369
rect 186502 700295 186558 700304
rect 135902 699816 135958 699825
rect 135902 699751 135958 699760
rect 137834 699816 137890 699825
rect 137834 699751 137890 699760
rect 135916 690713 135944 699751
rect 129922 690704 129978 690713
rect 129922 690639 129978 690648
rect 135902 690704 135958 690713
rect 135902 690639 135958 690648
rect 129936 686905 129964 690639
rect 129002 686896 129058 686905
rect 129002 686831 129058 686840
rect 129922 686896 129978 686905
rect 129922 686831 129978 686840
rect 129016 681873 129044 686831
rect 129002 681864 129058 681873
rect 129002 681799 129058 681808
rect 124862 681728 124918 681737
rect 124862 681663 124918 681672
rect 124876 670721 124904 681663
rect 123482 670712 123538 670721
rect 123482 670647 123538 670656
rect 124862 670712 124918 670721
rect 124862 670647 124918 670656
rect 123496 659569 123524 670647
rect 122102 659560 122158 659569
rect 122102 659495 122158 659504
rect 123482 659560 123538 659569
rect 123482 659495 123538 659504
rect 122116 650049 122144 659495
rect 120722 650040 120778 650049
rect 120722 649975 120778 649984
rect 122102 650040 122158 650049
rect 122102 649975 122158 649984
rect 120736 637537 120764 649975
rect 580262 644056 580318 644065
rect 580262 643991 580318 644000
rect 118790 637528 118846 637537
rect 118790 637463 118846 637472
rect 120722 637528 120778 637537
rect 120722 637463 120778 637472
rect 118804 634814 118832 637463
rect 118620 634786 118832 634814
rect 118620 630737 118648 634786
rect 116122 630728 116178 630737
rect 116122 630663 116178 630672
rect 118606 630728 118662 630737
rect 118606 630663 118662 630672
rect 116136 627881 116164 630663
rect 115202 627872 115258 627881
rect 115202 627807 115258 627816
rect 116122 627872 116178 627881
rect 116122 627807 116178 627816
rect 115216 612649 115244 627807
rect 111798 612640 111854 612649
rect 111798 612575 111854 612584
rect 115202 612640 115258 612649
rect 115202 612575 115258 612584
rect 111812 607889 111840 612575
rect 101402 607880 101458 607889
rect 101402 607815 101458 607824
rect 111798 607880 111854 607889
rect 111798 607815 111854 607824
rect 101416 597553 101444 607815
rect 98182 597544 98238 597553
rect 98182 597479 98238 597488
rect 101402 597544 101458 597553
rect 101402 597479 101458 597488
rect 98196 589529 98224 597479
rect 96618 589520 96674 589529
rect 96618 589455 96674 589464
rect 98182 589520 98238 589529
rect 98182 589455 98238 589464
rect 96632 588010 96660 589455
rect 96540 587982 96660 588010
rect 96540 586809 96568 587982
rect 96526 586800 96582 586809
rect 96526 586735 96582 586744
rect 89626 586392 89682 586401
rect 89626 586327 89682 586336
rect 89640 580961 89668 586327
rect 87602 580952 87658 580961
rect 87602 580887 87658 580896
rect 89626 580952 89682 580961
rect 89626 580887 89682 580896
rect 87616 575521 87644 580887
rect 84842 575512 84898 575521
rect 84842 575447 84898 575456
rect 87602 575512 87658 575521
rect 87602 575447 87658 575456
rect 84856 561649 84884 575447
rect 81438 561640 81494 561649
rect 81438 561575 81494 561584
rect 84842 561640 84898 561649
rect 84842 561575 84898 561584
rect 81452 559609 81480 561575
rect 76562 559600 76618 559609
rect 76562 559535 76618 559544
rect 81438 559600 81494 559609
rect 81438 559535 81494 559544
rect 76576 550633 76604 559535
rect 74630 550624 74686 550633
rect 74630 550559 74686 550568
rect 76562 550624 76618 550633
rect 76562 550559 76618 550568
rect 74644 545057 74672 550559
rect 73802 545048 73858 545057
rect 73802 544983 73858 544992
rect 74630 545048 74686 545057
rect 74630 544983 74686 544992
rect 73816 531321 73844 544983
rect 73802 531312 73858 531321
rect 73802 531247 73858 531256
rect 580078 484664 580134 484673
rect 580078 484599 580134 484608
rect 579894 431624 579950 431633
rect 579894 431559 579950 431568
rect 62762 409184 62818 409193
rect 62762 409119 62818 409128
rect 72974 409184 73030 409193
rect 72974 409119 73030 409128
rect 28998 408912 29054 408921
rect 28998 408847 29054 408856
rect 31758 408912 31814 408921
rect 31758 408847 31814 408856
rect 29012 407130 29040 408847
rect 28920 407102 29040 407130
rect 28920 406745 28948 407102
rect 25502 406736 25558 406745
rect 25502 406671 25558 406680
rect 28906 406736 28962 406745
rect 28906 406671 28962 406680
rect 25516 390697 25544 406671
rect 24122 390688 24178 390697
rect 24122 390623 24178 390632
rect 25502 390688 25558 390697
rect 25502 390623 25558 390632
rect 24136 380769 24164 390623
rect 22098 380760 22154 380769
rect 22098 380695 22154 380704
rect 24122 380760 24178 380769
rect 24122 380695 24178 380704
rect 22112 378185 22140 380695
rect 22098 378176 22154 378185
rect 22098 378111 22154 378120
rect 15842 377768 15898 377777
rect 15842 377703 15898 377712
rect 15856 371385 15884 377703
rect 62776 371385 62804 409119
rect 579710 378448 579766 378457
rect 579710 378383 579766 378392
rect 12346 371376 12402 371385
rect 12346 371311 12402 371320
rect 15842 371376 15898 371385
rect 15842 371311 15898 371320
rect 61382 371376 61438 371385
rect 61382 371311 61438 371320
rect 62762 371376 62818 371385
rect 62762 371311 62818 371320
rect 12254 143440 12310 143449
rect 12254 143375 12310 143384
rect 12360 4049 12388 371311
rect 61396 360233 61424 371311
rect 61382 360224 61438 360233
rect 61382 360159 61438 360168
rect 29642 359408 29698 359417
rect 29642 359343 29698 359352
rect 29656 324465 29684 359343
rect 26422 324456 26478 324465
rect 26344 324414 26422 324442
rect 26344 322946 26372 324414
rect 26422 324391 26478 324400
rect 29642 324456 29698 324465
rect 29642 324391 29698 324400
rect 26160 322918 26372 322946
rect 26160 321609 26188 322918
rect 22742 321600 22798 321609
rect 22742 321535 22798 321544
rect 26146 321600 26202 321609
rect 26146 321535 26202 321544
rect 22756 311953 22784 321535
rect 19982 311944 20038 311953
rect 19982 311879 20038 311888
rect 22742 311944 22798 311953
rect 22742 311879 22798 311888
rect 19996 304201 20024 311879
rect 17866 304192 17922 304201
rect 17866 304127 17922 304136
rect 19982 304192 20038 304201
rect 19982 304127 20038 304136
rect 17880 301889 17908 304127
rect 14462 301880 14518 301889
rect 14462 301815 14518 301824
rect 17866 301880 17922 301889
rect 17866 301815 17922 301824
rect 14476 284345 14504 301815
rect 12438 284336 12494 284345
rect 12438 284271 12494 284280
rect 14462 284336 14518 284345
rect 14462 284271 14518 284280
rect 12452 281489 12480 284271
rect 12438 281480 12494 281489
rect 12438 281415 12494 281424
rect 12346 4040 12402 4049
rect 12346 3975 12402 3984
rect 15198 4040 15254 4049
rect 15198 3975 15254 3984
rect 12162 3360 12218 3369
rect 12162 3295 12218 3304
rect 8114 1184 8170 1193
rect 8114 1119 8170 1128
rect 15212 1057 15240 3975
rect 21896 3046 22048 3074
rect 15198 1048 15254 1057
rect 15198 983 15254 992
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22020 377 22048 3046
rect 40420 3046 40480 3074
rect 59064 3046 59308 3074
rect 77648 3046 77984 3074
rect 96232 3046 96568 3074
rect 114816 3046 115152 3074
rect 40420 513 40448 3046
rect 59280 649 59308 3046
rect 77956 1329 77984 3046
rect 77942 1320 77998 1329
rect 77942 1255 77998 1264
rect 96540 921 96568 3046
rect 115124 1358 115152 3046
rect 133064 3046 133400 3074
rect 151832 3046 151984 3074
rect 170232 3046 170568 3074
rect 189152 3046 189488 3074
rect 207736 3046 208072 3074
rect 115112 1352 115164 1358
rect 115112 1294 115164 1300
rect 133064 1057 133092 3046
rect 151832 2689 151860 3046
rect 151818 2680 151874 2689
rect 151818 2615 151874 2624
rect 170232 1193 170260 3046
rect 189460 1193 189488 3046
rect 170218 1184 170274 1193
rect 170218 1119 170274 1128
rect 189446 1184 189502 1193
rect 189446 1119 189502 1128
rect 208044 1057 208072 3046
rect 226260 3046 226320 3074
rect 244904 3046 245240 3074
rect 133050 1048 133106 1057
rect 133050 983 133106 992
rect 208030 1048 208086 1057
rect 208030 983 208086 992
rect 226260 921 226288 3046
rect 244278 1320 244334 1329
rect 244278 1255 244280 1264
rect 244332 1255 244334 1264
rect 244280 1226 244332 1232
rect 96526 912 96582 921
rect 96526 847 96582 856
rect 224958 912 225014 921
rect 224958 847 225014 856
rect 226246 912 226302 921
rect 226246 847 226302 856
rect 224972 678 225000 847
rect 245212 785 245240 3046
rect 263428 3046 263488 3074
rect 282072 3046 282408 3074
rect 262864 1216 262916 1222
rect 262864 1158 262916 1164
rect 245198 776 245254 785
rect 245198 711 245254 720
rect 224960 672 225012 678
rect 59266 640 59322 649
rect 262876 649 262904 1158
rect 263428 649 263456 3046
rect 282184 1148 282236 1154
rect 282184 1090 282236 1096
rect 224960 614 225012 620
rect 262862 640 262918 649
rect 59266 575 59322 584
rect 262862 575 262918 584
rect 263414 640 263470 649
rect 263414 575 263470 584
rect 282196 513 282224 1090
rect 40406 504 40462 513
rect 22006 368 22062 377
rect 22006 303 22062 312
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 282182 504 282238 513
rect 40406 439 40462 448
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 282182 439 282238 448
rect 282380 105 282408 3046
rect 579620 1352 579672 1358
rect 579618 1320 579620 1329
rect 579672 1320 579674 1329
rect 579618 1255 579674 1264
rect 579724 1193 579752 378383
rect 579710 1184 579766 1193
rect 579710 1119 579766 1128
rect 579908 1057 579936 431559
rect 579894 1048 579950 1057
rect 579894 983 579950 992
rect 580092 921 580120 484599
rect 580078 912 580134 921
rect 580078 847 580134 856
rect 282366 96 282422 105
rect 282366 31 282422 40
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580276 105 580304 643991
rect 580446 591016 580502 591025
rect 580446 590951 580502 590960
rect 580354 511320 580410 511329
rect 580354 511255 580410 511264
rect 580368 1290 580396 511255
rect 580356 1284 580408 1290
rect 580356 1226 580408 1232
rect 580354 912 580410 921
rect 580354 847 580410 856
rect 580368 678 580396 847
rect 580356 672 580408 678
rect 580460 649 580488 590951
rect 580906 537840 580962 537849
rect 580906 537775 580962 537784
rect 580538 458144 580594 458153
rect 580538 458079 580594 458088
rect 580552 1222 580580 458079
rect 580630 404968 580686 404977
rect 580630 404903 580686 404912
rect 580540 1216 580592 1222
rect 580540 1158 580592 1164
rect 580644 1154 580672 404903
rect 580722 351928 580778 351937
rect 580722 351863 580778 351872
rect 580632 1148 580684 1154
rect 580632 1090 580684 1096
rect 580356 614 580408 620
rect 580446 640 580502 649
rect 580446 575 580502 584
rect 580736 377 580764 351863
rect 580920 785 580948 537775
rect 580906 776 580962 785
rect 580906 711 580962 720
rect 580722 368 580778 377
rect 580722 303 580778 312
rect 580262 96 580318 105
rect 580262 31 580318 40
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 12070 700576 12126 700632
rect 56782 700576 56838 700632
rect 9586 700304 9642 700360
rect 9586 236136 9642 236192
rect 12254 700440 12310 700496
rect 12162 281424 12218 281480
rect 12070 49816 12126 49872
rect 71778 531256 71834 531312
rect 66902 522960 66958 523016
rect 71686 522960 71742 523016
rect 65522 506504 65578 506560
rect 66902 506504 66958 506560
rect 65522 487328 65578 487384
rect 62762 487056 62818 487112
rect 60738 475360 60794 475416
rect 62762 475360 62818 475416
rect 58622 473184 58678 473240
rect 60646 473184 60702 473240
rect 56874 459584 56930 459640
rect 58622 459584 58678 459640
rect 54482 458224 54538 458280
rect 56874 458224 56930 458280
rect 53102 446392 53158 446448
rect 54482 446392 54538 446448
rect 53102 434696 53158 434752
rect 46938 434560 46994 434616
rect 42798 422320 42854 422376
rect 46846 422320 46902 422376
rect 38566 418240 38622 418296
rect 42706 418240 42762 418296
rect 38566 412664 38622 412720
rect 31758 412528 31814 412584
rect 121642 700440 121698 700496
rect 186502 700304 186558 700360
rect 135902 699760 135958 699816
rect 137834 699760 137890 699816
rect 129922 690648 129978 690704
rect 135902 690648 135958 690704
rect 129002 686840 129058 686896
rect 129922 686840 129978 686896
rect 129002 681808 129058 681864
rect 124862 681672 124918 681728
rect 123482 670656 123538 670712
rect 124862 670656 124918 670712
rect 122102 659504 122158 659560
rect 123482 659504 123538 659560
rect 120722 649984 120778 650040
rect 122102 649984 122158 650040
rect 580262 644000 580318 644056
rect 118790 637472 118846 637528
rect 120722 637472 120778 637528
rect 116122 630672 116178 630728
rect 118606 630672 118662 630728
rect 115202 627816 115258 627872
rect 116122 627816 116178 627872
rect 111798 612584 111854 612640
rect 115202 612584 115258 612640
rect 101402 607824 101458 607880
rect 111798 607824 111854 607880
rect 98182 597488 98238 597544
rect 101402 597488 101458 597544
rect 96618 589464 96674 589520
rect 98182 589464 98238 589520
rect 96526 586744 96582 586800
rect 89626 586336 89682 586392
rect 87602 580896 87658 580952
rect 89626 580896 89682 580952
rect 84842 575456 84898 575512
rect 87602 575456 87658 575512
rect 81438 561584 81494 561640
rect 84842 561584 84898 561640
rect 76562 559544 76618 559600
rect 81438 559544 81494 559600
rect 74630 550568 74686 550624
rect 76562 550568 76618 550624
rect 73802 544992 73858 545048
rect 74630 544992 74686 545048
rect 73802 531256 73858 531312
rect 580078 484608 580134 484664
rect 579894 431568 579950 431624
rect 62762 409128 62818 409184
rect 72974 409128 73030 409184
rect 28998 408856 29054 408912
rect 31758 408856 31814 408912
rect 25502 406680 25558 406736
rect 28906 406680 28962 406736
rect 24122 390632 24178 390688
rect 25502 390632 25558 390688
rect 22098 380704 22154 380760
rect 24122 380704 24178 380760
rect 22098 378120 22154 378176
rect 15842 377712 15898 377768
rect 579710 378392 579766 378448
rect 12346 371320 12402 371376
rect 15842 371320 15898 371376
rect 61382 371320 61438 371376
rect 62762 371320 62818 371376
rect 12254 143384 12310 143440
rect 61382 360168 61438 360224
rect 29642 359352 29698 359408
rect 26422 324400 26478 324456
rect 29642 324400 29698 324456
rect 22742 321544 22798 321600
rect 26146 321544 26202 321600
rect 19982 311888 20038 311944
rect 22742 311888 22798 311944
rect 17866 304136 17922 304192
rect 19982 304136 20038 304192
rect 14462 301824 14518 301880
rect 17866 301824 17922 301880
rect 12438 284280 12494 284336
rect 14462 284280 14518 284336
rect 12438 281424 12494 281480
rect 12346 3984 12402 4040
rect 15198 3984 15254 4040
rect 12162 3304 12218 3360
rect 8114 1128 8170 1184
rect 15198 992 15254 1048
rect 77942 1264 77998 1320
rect 151818 2624 151874 2680
rect 170218 1128 170274 1184
rect 189446 1128 189502 1184
rect 133050 992 133106 1048
rect 208030 992 208086 1048
rect 244278 1284 244334 1320
rect 244278 1264 244280 1284
rect 244280 1264 244332 1284
rect 244332 1264 244334 1284
rect 96526 856 96582 912
rect 224958 856 225014 912
rect 226246 856 226302 912
rect 245198 720 245254 776
rect 59266 584 59322 640
rect 262862 584 262918 640
rect 263414 584 263470 640
rect 22006 312 22062 368
rect 40406 448 40462 504
rect 282182 448 282238 504
rect 579618 1300 579620 1320
rect 579620 1300 579672 1320
rect 579672 1300 579674 1320
rect 579618 1264 579674 1300
rect 579710 1128 579766 1184
rect 579894 992 579950 1048
rect 580078 856 580134 912
rect 282366 40 282422 96
rect 580446 590960 580502 591016
rect 580354 511264 580410 511320
rect 580354 856 580410 912
rect 580906 537784 580962 537840
rect 580538 458088 580594 458144
rect 580630 404912 580686 404968
rect 580722 351872 580778 351928
rect 580446 584 580502 640
rect 580906 720 580962 776
rect 580722 312 580778 368
rect 580262 40 580318 96
<< metal3 >>
rect 12065 700634 12131 700637
rect 56777 700634 56843 700637
rect 12065 700632 56843 700634
rect 12065 700576 12070 700632
rect 12126 700576 56782 700632
rect 56838 700576 56843 700632
rect 12065 700574 56843 700576
rect 12065 700571 12131 700574
rect 56777 700571 56843 700574
rect 12249 700498 12315 700501
rect 121637 700498 121703 700501
rect 12249 700496 121703 700498
rect 12249 700440 12254 700496
rect 12310 700440 121642 700496
rect 121698 700440 121703 700496
rect 12249 700438 121703 700440
rect 12249 700435 12315 700438
rect 121637 700435 121703 700438
rect 9581 700362 9647 700365
rect 186497 700362 186563 700365
rect 9581 700360 186563 700362
rect 9581 700304 9586 700360
rect 9642 700304 186502 700360
rect 186558 700304 186563 700360
rect 9581 700302 186563 700304
rect 9581 700299 9647 700302
rect 186497 700299 186563 700302
rect 135897 699818 135963 699821
rect 137829 699818 137895 699821
rect 135897 699816 137895 699818
rect 135897 699760 135902 699816
rect 135958 699760 137834 699816
rect 137890 699760 137895 699816
rect 135897 699758 137895 699760
rect 135897 699755 135963 699758
rect 137829 699755 137895 699758
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect 129917 690706 129983 690709
rect 135897 690706 135963 690709
rect 129917 690704 135963 690706
rect 129917 690648 129922 690704
rect 129978 690648 135902 690704
rect 135958 690648 135963 690704
rect 129917 690646 135963 690648
rect 129917 690643 129983 690646
rect 135897 690643 135963 690646
rect 128997 686898 129063 686901
rect 129917 686898 129983 686901
rect 128997 686896 129983 686898
rect 128997 686840 129002 686896
rect 129058 686840 129922 686896
rect 129978 686840 129983 686896
rect 128997 686838 129983 686840
rect 128997 686835 129063 686838
rect 129917 686835 129983 686838
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect 128997 681866 129063 681869
rect 127022 681864 129063 681866
rect 127022 681808 129002 681864
rect 129058 681808 129063 681864
rect 127022 681806 129063 681808
rect 124857 681730 124923 681733
rect 127022 681730 127082 681806
rect 128997 681803 129063 681806
rect 124857 681728 127082 681730
rect 124857 681672 124862 681728
rect 124918 681672 127082 681728
rect 124857 681670 127082 681672
rect 124857 681667 124923 681670
rect -960 671108 480 671348
rect 123477 670714 123543 670717
rect 124857 670714 124923 670717
rect 123477 670712 124923 670714
rect 123477 670656 123482 670712
rect 123538 670656 124862 670712
rect 124918 670656 124923 670712
rect 123477 670654 124923 670656
rect 123477 670651 123543 670654
rect 124857 670651 124923 670654
rect 583520 670564 584960 670804
rect 122097 659562 122163 659565
rect 123477 659562 123543 659565
rect 122097 659560 123543 659562
rect 122097 659504 122102 659560
rect 122158 659504 123482 659560
rect 123538 659504 123543 659560
rect 122097 659502 123543 659504
rect 122097 659499 122163 659502
rect 123477 659499 123543 659502
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect 120717 650042 120783 650045
rect 122097 650042 122163 650045
rect 120717 650040 122163 650042
rect 120717 649984 120722 650040
rect 120778 649984 122102 650040
rect 122158 649984 122163 650040
rect 120717 649982 122163 649984
rect 120717 649979 120783 649982
rect 122097 649979 122163 649982
rect -960 644996 480 645236
rect 580257 644058 580323 644061
rect 583520 644058 584960 644148
rect 580257 644056 584960 644058
rect 580257 644000 580262 644056
rect 580318 644000 584960 644056
rect 580257 643998 584960 644000
rect 580257 643995 580323 643998
rect 583520 643908 584960 643998
rect 118785 637530 118851 637533
rect 120717 637530 120783 637533
rect 118785 637528 120783 637530
rect 118785 637472 118790 637528
rect 118846 637472 120722 637528
rect 120778 637472 120783 637528
rect 118785 637470 120783 637472
rect 118785 637467 118851 637470
rect 120717 637467 120783 637470
rect -960 631940 480 632180
rect 116117 630730 116183 630733
rect 118601 630730 118667 630733
rect 116117 630728 118667 630730
rect 116117 630672 116122 630728
rect 116178 630672 118606 630728
rect 118662 630672 118667 630728
rect 583520 630716 584960 630956
rect 116117 630670 118667 630672
rect 116117 630667 116183 630670
rect 118601 630667 118667 630670
rect 115197 627874 115263 627877
rect 116117 627874 116183 627877
rect 115197 627872 116183 627874
rect 115197 627816 115202 627872
rect 115258 627816 116122 627872
rect 116178 627816 116183 627872
rect 115197 627814 116183 627816
rect 115197 627811 115263 627814
rect 116117 627811 116183 627814
rect -960 619020 480 619260
rect 580390 617476 580396 617540
rect 580460 617538 580466 617540
rect 583520 617538 584960 617628
rect 580460 617478 584960 617538
rect 580460 617476 580466 617478
rect 583520 617388 584960 617478
rect 111793 612642 111859 612645
rect 115197 612642 115263 612645
rect 111793 612640 115263 612642
rect 111793 612584 111798 612640
rect 111854 612584 115202 612640
rect 115258 612584 115263 612640
rect 111793 612582 115263 612584
rect 111793 612579 111859 612582
rect 115197 612579 115263 612582
rect 101397 607882 101463 607885
rect 111793 607882 111859 607885
rect 101397 607880 111859 607882
rect 101397 607824 101402 607880
rect 101458 607824 111798 607880
rect 111854 607824 111859 607880
rect 101397 607822 111859 607824
rect 101397 607819 101463 607822
rect 111793 607819 111859 607822
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect 98177 597546 98243 597549
rect 101397 597546 101463 597549
rect 98177 597544 101463 597546
rect 98177 597488 98182 597544
rect 98238 597488 101402 597544
rect 101458 597488 101463 597544
rect 98177 597486 101463 597488
rect 98177 597483 98243 597486
rect 101397 597483 101463 597486
rect -960 592908 480 593148
rect 580441 591018 580507 591021
rect 583520 591018 584960 591108
rect 580441 591016 584960 591018
rect 580441 590960 580446 591016
rect 580502 590960 584960 591016
rect 580441 590958 584960 590960
rect 580441 590955 580507 590958
rect 583520 590868 584960 590958
rect 96613 589522 96679 589525
rect 98177 589522 98243 589525
rect 96613 589520 98243 589522
rect 96613 589464 96618 589520
rect 96674 589464 98182 589520
rect 98238 589464 98243 589520
rect 96613 589462 98243 589464
rect 96613 589459 96679 589462
rect 98177 589459 98243 589462
rect 96521 586802 96587 586805
rect 95190 586800 96587 586802
rect 95190 586744 96526 586800
rect 96582 586744 96587 586800
rect 95190 586742 96587 586744
rect 89621 586394 89687 586397
rect 95190 586394 95250 586742
rect 96521 586739 96587 586742
rect 89621 586392 95250 586394
rect 89621 586336 89626 586392
rect 89682 586336 95250 586392
rect 89621 586334 95250 586336
rect 89621 586331 89687 586334
rect 87597 580954 87663 580957
rect 89621 580954 89687 580957
rect 87597 580952 89687 580954
rect 87597 580896 87602 580952
rect 87658 580896 89626 580952
rect 89682 580896 89687 580952
rect 87597 580894 89687 580896
rect 87597 580891 87663 580894
rect 89621 580891 89687 580894
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect 84837 575514 84903 575517
rect 87597 575514 87663 575517
rect 84837 575512 87663 575514
rect 84837 575456 84842 575512
rect 84898 575456 87602 575512
rect 87658 575456 87663 575512
rect 84837 575454 87663 575456
rect 84837 575451 84903 575454
rect 87597 575451 87663 575454
rect -960 566796 480 567036
rect 580574 564300 580580 564364
rect 580644 564362 580650 564364
rect 583520 564362 584960 564452
rect 580644 564302 584960 564362
rect 580644 564300 580650 564302
rect 583520 564212 584960 564302
rect 81433 561642 81499 561645
rect 84837 561642 84903 561645
rect 81433 561640 84903 561642
rect 81433 561584 81438 561640
rect 81494 561584 84842 561640
rect 84898 561584 84903 561640
rect 81433 561582 84903 561584
rect 81433 561579 81499 561582
rect 84837 561579 84903 561582
rect 76557 559602 76623 559605
rect 81433 559602 81499 559605
rect 76557 559600 81499 559602
rect 76557 559544 76562 559600
rect 76618 559544 81438 559600
rect 81494 559544 81499 559600
rect 76557 559542 81499 559544
rect 76557 559539 76623 559542
rect 81433 559539 81499 559542
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect 74625 550626 74691 550629
rect 76557 550626 76623 550629
rect 74625 550624 76623 550626
rect 74625 550568 74630 550624
rect 74686 550568 76562 550624
rect 76618 550568 76623 550624
rect 74625 550566 76623 550568
rect 74625 550563 74691 550566
rect 76557 550563 76623 550566
rect 73797 545050 73863 545053
rect 74625 545050 74691 545053
rect 73797 545048 74691 545050
rect 73797 544992 73802 545048
rect 73858 544992 74630 545048
rect 74686 544992 74691 545048
rect 73797 544990 74691 544992
rect 73797 544987 73863 544990
rect 74625 544987 74691 544990
rect -960 540684 480 540924
rect 580901 537842 580967 537845
rect 583520 537842 584960 537932
rect 580901 537840 584960 537842
rect 580901 537784 580906 537840
rect 580962 537784 584960 537840
rect 580901 537782 584960 537784
rect 580901 537779 580967 537782
rect 583520 537692 584960 537782
rect 71773 531314 71839 531317
rect 73797 531314 73863 531317
rect 71773 531312 73863 531314
rect 71773 531256 71778 531312
rect 71834 531256 73802 531312
rect 73858 531256 73863 531312
rect 71773 531254 73863 531256
rect 71773 531251 71839 531254
rect 73797 531251 73863 531254
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect 66897 523018 66963 523021
rect 71681 523018 71747 523021
rect 66897 523016 71747 523018
rect 66897 522960 66902 523016
rect 66958 522960 71686 523016
rect 71742 522960 71747 523016
rect 66897 522958 71747 522960
rect 66897 522955 66963 522958
rect 71681 522955 71747 522958
rect -960 514708 480 514948
rect 580349 511322 580415 511325
rect 583520 511322 584960 511412
rect 580349 511320 584960 511322
rect 580349 511264 580354 511320
rect 580410 511264 584960 511320
rect 580349 511262 584960 511264
rect 580349 511259 580415 511262
rect 583520 511172 584960 511262
rect 65517 506562 65583 506565
rect 66897 506562 66963 506565
rect 65517 506560 66963 506562
rect 65517 506504 65522 506560
rect 65578 506504 66902 506560
rect 66958 506504 66963 506560
rect 65517 506502 66963 506504
rect 65517 506499 65583 506502
rect 66897 506499 66963 506502
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 65517 487386 65583 487389
rect 64830 487384 65583 487386
rect 64830 487328 65522 487384
rect 65578 487328 65583 487384
rect 64830 487326 65583 487328
rect 62757 487114 62823 487117
rect 64830 487114 64890 487326
rect 65517 487323 65583 487326
rect 62757 487112 64890 487114
rect 62757 487056 62762 487112
rect 62818 487056 64890 487112
rect 62757 487054 64890 487056
rect 62757 487051 62823 487054
rect 580073 484666 580139 484669
rect 583520 484666 584960 484756
rect 580073 484664 584960 484666
rect 580073 484608 580078 484664
rect 580134 484608 584960 484664
rect 580073 484606 584960 484608
rect 580073 484603 580139 484606
rect 583520 484516 584960 484606
rect -960 475540 480 475780
rect 60733 475418 60799 475421
rect 62757 475418 62823 475421
rect 60733 475416 62823 475418
rect 60733 475360 60738 475416
rect 60794 475360 62762 475416
rect 62818 475360 62823 475416
rect 60733 475358 62823 475360
rect 60733 475355 60799 475358
rect 62757 475355 62823 475358
rect 58617 473242 58683 473245
rect 60641 473242 60707 473245
rect 58617 473240 60707 473242
rect 58617 473184 58622 473240
rect 58678 473184 60646 473240
rect 60702 473184 60707 473240
rect 58617 473182 60707 473184
rect 58617 473179 58683 473182
rect 60641 473179 60707 473182
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 56869 459642 56935 459645
rect 58617 459642 58683 459645
rect 56869 459640 58683 459642
rect 56869 459584 56874 459640
rect 56930 459584 58622 459640
rect 58678 459584 58683 459640
rect 56869 459582 58683 459584
rect 56869 459579 56935 459582
rect 58617 459579 58683 459582
rect 54477 458282 54543 458285
rect 56869 458282 56935 458285
rect 54477 458280 56935 458282
rect 54477 458224 54482 458280
rect 54538 458224 56874 458280
rect 56930 458224 56935 458280
rect 54477 458222 56935 458224
rect 54477 458219 54543 458222
rect 56869 458219 56935 458222
rect 580533 458146 580599 458149
rect 583520 458146 584960 458236
rect 580533 458144 584960 458146
rect 580533 458088 580538 458144
rect 580594 458088 584960 458144
rect 580533 458086 584960 458088
rect 580533 458083 580599 458086
rect 583520 457996 584960 458086
rect -960 449428 480 449668
rect 53097 446450 53163 446453
rect 54477 446450 54543 446453
rect 53097 446448 54543 446450
rect 53097 446392 53102 446448
rect 53158 446392 54482 446448
rect 54538 446392 54543 446448
rect 53097 446390 54543 446392
rect 53097 446387 53163 446390
rect 54477 446387 54543 446390
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 53097 434754 53163 434757
rect 51030 434752 53163 434754
rect 51030 434696 53102 434752
rect 53158 434696 53163 434752
rect 51030 434694 53163 434696
rect 46933 434618 46999 434621
rect 51030 434618 51090 434694
rect 53097 434691 53163 434694
rect 46933 434616 51090 434618
rect 46933 434560 46938 434616
rect 46994 434560 51090 434616
rect 46933 434558 51090 434560
rect 46933 434555 46999 434558
rect 579889 431626 579955 431629
rect 583520 431626 584960 431716
rect 579889 431624 584960 431626
rect 579889 431568 579894 431624
rect 579950 431568 584960 431624
rect 579889 431566 584960 431568
rect 579889 431563 579955 431566
rect 583520 431476 584960 431566
rect -960 423452 480 423692
rect 42793 422378 42859 422381
rect 46841 422378 46907 422381
rect 42793 422376 46907 422378
rect 42793 422320 42798 422376
rect 42854 422320 46846 422376
rect 46902 422320 46907 422376
rect 42793 422318 46907 422320
rect 42793 422315 42859 422318
rect 46841 422315 46907 422318
rect 38561 418298 38627 418301
rect 42701 418298 42767 418301
rect 38561 418296 42767 418298
rect 38561 418240 38566 418296
rect 38622 418240 42706 418296
rect 42762 418240 42767 418296
rect 38561 418238 42767 418240
rect 38561 418235 38627 418238
rect 42701 418235 42767 418238
rect 583520 418148 584960 418388
rect 38561 412722 38627 412725
rect 34470 412720 38627 412722
rect 34470 412664 38566 412720
rect 38622 412664 38627 412720
rect 34470 412662 38627 412664
rect 31753 412586 31819 412589
rect 34470 412586 34530 412662
rect 38561 412659 38627 412662
rect 31753 412584 34530 412586
rect 31753 412528 31758 412584
rect 31814 412528 34530 412584
rect 31753 412526 34530 412528
rect 31753 412523 31819 412526
rect -960 410396 480 410636
rect 62757 409186 62823 409189
rect 72969 409186 73035 409189
rect 62757 409184 73035 409186
rect 62757 409128 62762 409184
rect 62818 409128 72974 409184
rect 73030 409128 73035 409184
rect 62757 409126 73035 409128
rect 62757 409123 62823 409126
rect 72969 409123 73035 409126
rect 28993 408914 29059 408917
rect 31753 408914 31819 408917
rect 28993 408912 31819 408914
rect 28993 408856 28998 408912
rect 29054 408856 31758 408912
rect 31814 408856 31819 408912
rect 28993 408854 31819 408856
rect 28993 408851 29059 408854
rect 31753 408851 31819 408854
rect 25497 406738 25563 406741
rect 28901 406738 28967 406741
rect 25497 406736 28967 406738
rect 25497 406680 25502 406736
rect 25558 406680 28906 406736
rect 28962 406680 28967 406736
rect 25497 406678 28967 406680
rect 25497 406675 25563 406678
rect 28901 406675 28967 406678
rect 580625 404970 580691 404973
rect 583520 404970 584960 405060
rect 580625 404968 584960 404970
rect 580625 404912 580630 404968
rect 580686 404912 584960 404968
rect 580625 404910 584960 404912
rect 580625 404907 580691 404910
rect 583520 404820 584960 404910
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect 24117 390690 24183 390693
rect 25497 390690 25563 390693
rect 24117 390688 25563 390690
rect 24117 390632 24122 390688
rect 24178 390632 25502 390688
rect 25558 390632 25563 390688
rect 24117 390630 25563 390632
rect 24117 390627 24183 390630
rect 25497 390627 25563 390630
rect -960 384284 480 384524
rect 22093 380762 22159 380765
rect 24117 380762 24183 380765
rect 22093 380760 24183 380762
rect 22093 380704 22098 380760
rect 22154 380704 24122 380760
rect 24178 380704 24183 380760
rect 22093 380702 24183 380704
rect 22093 380699 22159 380702
rect 24117 380699 24183 380702
rect 579705 378450 579771 378453
rect 583520 378450 584960 378540
rect 579705 378448 584960 378450
rect 579705 378392 579710 378448
rect 579766 378392 584960 378448
rect 579705 378390 584960 378392
rect 579705 378387 579771 378390
rect 583520 378300 584960 378390
rect 22093 378178 22159 378181
rect 19198 378176 22159 378178
rect 19198 378120 22098 378176
rect 22154 378120 22159 378176
rect 19198 378118 22159 378120
rect 15837 377770 15903 377773
rect 19198 377770 19258 378118
rect 22093 378115 22159 378118
rect 15837 377768 19258 377770
rect 15837 377712 15842 377768
rect 15898 377712 19258 377768
rect 15837 377710 19258 377712
rect 15837 377707 15903 377710
rect -960 371228 480 371468
rect 12341 371378 12407 371381
rect 15837 371378 15903 371381
rect 12341 371376 15903 371378
rect 12341 371320 12346 371376
rect 12402 371320 15842 371376
rect 15898 371320 15903 371376
rect 12341 371318 15903 371320
rect 12341 371315 12407 371318
rect 15837 371315 15903 371318
rect 61377 371378 61443 371381
rect 62757 371378 62823 371381
rect 61377 371376 62823 371378
rect 61377 371320 61382 371376
rect 61438 371320 62762 371376
rect 62818 371320 62823 371376
rect 61377 371318 62823 371320
rect 61377 371315 61443 371318
rect 62757 371315 62823 371318
rect 583520 364972 584960 365212
rect 61377 360226 61443 360229
rect 59310 360224 61443 360226
rect 59310 360168 61382 360224
rect 61438 360168 61443 360224
rect 59310 360166 61443 360168
rect 29637 359410 29703 359413
rect 59310 359410 59370 360166
rect 61377 360163 61443 360166
rect 29637 359408 59370 359410
rect 29637 359352 29642 359408
rect 29698 359352 59370 359408
rect 29637 359350 59370 359352
rect 29637 359347 29703 359350
rect -960 358308 480 358548
rect 580717 351930 580783 351933
rect 583520 351930 584960 352020
rect 580717 351928 584960 351930
rect 580717 351872 580722 351928
rect 580778 351872 584960 351928
rect 580717 351870 584960 351872
rect 580717 351867 580783 351870
rect 583520 351780 584960 351870
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect 26417 324458 26483 324461
rect 29637 324458 29703 324461
rect 26417 324456 29703 324458
rect 26417 324400 26422 324456
rect 26478 324400 29642 324456
rect 29698 324400 29703 324456
rect 26417 324398 29703 324400
rect 26417 324395 26483 324398
rect 29637 324395 29703 324398
rect 22737 321602 22803 321605
rect 26141 321602 26207 321605
rect 22737 321600 26207 321602
rect 22737 321544 22742 321600
rect 22798 321544 26146 321600
rect 26202 321544 26207 321600
rect 22737 321542 26207 321544
rect 22737 321539 22803 321542
rect 26141 321539 26207 321542
rect -960 319140 480 319380
rect 19977 311946 20043 311949
rect 22737 311946 22803 311949
rect 19977 311944 22803 311946
rect 19977 311888 19982 311944
rect 20038 311888 22742 311944
rect 22798 311888 22803 311944
rect 583520 311932 584960 312172
rect 19977 311886 22803 311888
rect 19977 311883 20043 311886
rect 22737 311883 22803 311886
rect -960 306084 480 306324
rect 17861 304194 17927 304197
rect 19977 304194 20043 304197
rect 17861 304192 20043 304194
rect 17861 304136 17866 304192
rect 17922 304136 19982 304192
rect 20038 304136 20043 304192
rect 17861 304134 20043 304136
rect 17861 304131 17927 304134
rect 19977 304131 20043 304134
rect 14457 301882 14523 301885
rect 17861 301882 17927 301885
rect 14457 301880 17927 301882
rect 14457 301824 14462 301880
rect 14518 301824 17866 301880
rect 17922 301824 17927 301880
rect 14457 301822 17927 301824
rect 14457 301819 14523 301822
rect 17861 301819 17927 301822
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect 12433 284338 12499 284341
rect 14457 284338 14523 284341
rect 12433 284336 14523 284338
rect 12433 284280 12438 284336
rect 12494 284280 14462 284336
rect 14518 284280 14523 284336
rect 12433 284278 14523 284280
rect 12433 284275 12499 284278
rect 14457 284275 14523 284278
rect 12157 281482 12223 281485
rect 12433 281482 12499 281485
rect 12157 281480 12499 281482
rect 12157 281424 12162 281480
rect 12218 281424 12438 281480
rect 12494 281424 12499 281480
rect 12157 281422 12499 281424
rect 12157 281419 12223 281422
rect 12433 281419 12499 281422
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 9581 236194 9647 236197
rect 9581 236192 12052 236194
rect 9581 236136 9586 236192
rect 9642 236136 12052 236192
rect 9581 236134 12052 236136
rect 9581 236131 9647 236134
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 12249 143442 12315 143445
rect 12206 143440 12315 143442
rect 12206 143384 12254 143440
rect 12310 143384 12315 143440
rect 12206 143379 12315 143384
rect 12206 142868 12266 143379
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 12065 49874 12131 49877
rect 12022 49872 12131 49874
rect 12022 49816 12070 49872
rect 12126 49816 12131 49872
rect 12022 49811 12131 49816
rect 12022 49572 12082 49811
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
rect 12341 4042 12407 4045
rect 15193 4042 15259 4045
rect 12341 4040 15259 4042
rect 12341 3984 12346 4040
rect 12402 3984 15198 4040
rect 15254 3984 15259 4040
rect 12341 3982 15259 3984
rect 12341 3979 12407 3982
rect 15193 3979 15259 3982
rect 12157 3362 12223 3365
rect 12157 3360 31034 3362
rect 12157 3304 12162 3360
rect 12218 3304 31034 3360
rect 12157 3302 31034 3304
rect 12157 3299 12223 3302
rect 30974 2682 31034 3302
rect 151813 2682 151879 2685
rect 30974 2680 151879 2682
rect 30974 2624 151818 2680
rect 151874 2624 151879 2680
rect 30974 2622 151879 2624
rect 151813 2619 151879 2622
rect 77937 1322 78003 1325
rect 244273 1322 244339 1325
rect 77937 1320 244339 1322
rect 77937 1264 77942 1320
rect 77998 1264 244278 1320
rect 244334 1264 244339 1320
rect 77937 1262 244339 1264
rect 77937 1259 78003 1262
rect 244273 1259 244339 1262
rect 579613 1322 579679 1325
rect 580390 1322 580396 1324
rect 579613 1320 580396 1322
rect 579613 1264 579618 1320
rect 579674 1264 580396 1320
rect 579613 1262 580396 1264
rect 579613 1259 579679 1262
rect 580390 1260 580396 1262
rect 580460 1260 580466 1324
rect 8109 1186 8175 1189
rect 170213 1186 170279 1189
rect 8109 1184 170279 1186
rect 8109 1128 8114 1184
rect 8170 1128 170218 1184
rect 170274 1128 170279 1184
rect 8109 1126 170279 1128
rect 8109 1123 8175 1126
rect 170213 1123 170279 1126
rect 189441 1186 189507 1189
rect 579705 1186 579771 1189
rect 189441 1184 579771 1186
rect 189441 1128 189446 1184
rect 189502 1128 579710 1184
rect 579766 1128 579771 1184
rect 189441 1126 579771 1128
rect 189441 1123 189507 1126
rect 579705 1123 579771 1126
rect 15193 1050 15259 1053
rect 133045 1050 133111 1053
rect 15193 1048 133111 1050
rect 15193 992 15198 1048
rect 15254 992 133050 1048
rect 133106 992 133111 1048
rect 15193 990 133111 992
rect 15193 987 15259 990
rect 133045 987 133111 990
rect 208025 1050 208091 1053
rect 579889 1050 579955 1053
rect 208025 1048 579955 1050
rect 208025 992 208030 1048
rect 208086 992 579894 1048
rect 579950 992 579955 1048
rect 208025 990 579955 992
rect 208025 987 208091 990
rect 579889 987 579955 990
rect 96521 914 96587 917
rect 224953 914 225019 917
rect 96521 912 225019 914
rect 96521 856 96526 912
rect 96582 856 224958 912
rect 225014 856 225019 912
rect 96521 854 225019 856
rect 96521 851 96587 854
rect 224953 851 225019 854
rect 226241 914 226307 917
rect 580073 914 580139 917
rect 226241 912 580139 914
rect 226241 856 226246 912
rect 226302 856 580078 912
rect 580134 856 580139 912
rect 226241 854 580139 856
rect 226241 851 226307 854
rect 580073 851 580139 854
rect 580349 914 580415 917
rect 580574 914 580580 916
rect 580349 912 580580 914
rect 580349 856 580354 912
rect 580410 856 580580 912
rect 580349 854 580580 856
rect 580349 851 580415 854
rect 580574 852 580580 854
rect 580644 852 580650 916
rect 245193 778 245259 781
rect 580901 778 580967 781
rect 245193 776 580967 778
rect 245193 720 245198 776
rect 245254 720 580906 776
rect 580962 720 580967 776
rect 245193 718 580967 720
rect 245193 715 245259 718
rect 580901 715 580967 718
rect 59261 642 59327 645
rect 262857 642 262923 645
rect 59261 640 262923 642
rect 59261 584 59266 640
rect 59322 584 262862 640
rect 262918 584 262923 640
rect 59261 582 262923 584
rect 59261 579 59327 582
rect 262857 579 262923 582
rect 263409 642 263475 645
rect 580441 642 580507 645
rect 263409 640 580507 642
rect 263409 584 263414 640
rect 263470 584 580446 640
rect 580502 584 580507 640
rect 263409 582 580507 584
rect 263409 579 263475 582
rect 580441 579 580507 582
rect 40401 506 40467 509
rect 282177 506 282243 509
rect 40401 504 282243 506
rect 40401 448 40406 504
rect 40462 448 282182 504
rect 282238 448 282243 504
rect 40401 446 282243 448
rect 40401 443 40467 446
rect 282177 443 282243 446
rect 22001 370 22067 373
rect 580717 370 580783 373
rect 22001 368 580783 370
rect 22001 312 22006 368
rect 22062 312 580722 368
rect 580778 312 580783 368
rect 22001 310 580783 312
rect 22001 307 22067 310
rect 580717 307 580783 310
rect 282361 98 282427 101
rect 580257 98 580323 101
rect 282361 96 580323 98
rect 282361 40 282366 96
rect 282422 40 580262 96
rect 580318 40 580323 96
rect 282361 38 580323 40
rect 282361 35 282427 38
rect 580257 35 580323 38
<< via3 >>
rect 580396 617476 580460 617540
rect 580580 564300 580644 564364
rect 580396 1260 580460 1324
rect 580580 852 580644 916
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711002 -8694 711558
rect -8138 711002 -8106 711558
rect -8726 677494 -8106 711002
rect -8726 676938 -8694 677494
rect -8138 676938 -8106 677494
rect -8726 641494 -8106 676938
rect -8726 640938 -8694 641494
rect -8138 640938 -8106 641494
rect -8726 605494 -8106 640938
rect -8726 604938 -8694 605494
rect -8138 604938 -8106 605494
rect -8726 569494 -8106 604938
rect -8726 568938 -8694 569494
rect -8138 568938 -8106 569494
rect -8726 533494 -8106 568938
rect -8726 532938 -8694 533494
rect -8138 532938 -8106 533494
rect -8726 497494 -8106 532938
rect -8726 496938 -8694 497494
rect -8138 496938 -8106 497494
rect -8726 461494 -8106 496938
rect -8726 460938 -8694 461494
rect -8138 460938 -8106 461494
rect -8726 425494 -8106 460938
rect -8726 424938 -8694 425494
rect -8138 424938 -8106 425494
rect -8726 389494 -8106 424938
rect -8726 388938 -8694 389494
rect -8138 388938 -8106 389494
rect -8726 353494 -8106 388938
rect -8726 352938 -8694 353494
rect -8138 352938 -8106 353494
rect -8726 317494 -8106 352938
rect -8726 316938 -8694 317494
rect -8138 316938 -8106 317494
rect -8726 281494 -8106 316938
rect -8726 280938 -8694 281494
rect -8138 280938 -8106 281494
rect -8726 245494 -8106 280938
rect -8726 244938 -8694 245494
rect -8138 244938 -8106 245494
rect -8726 209494 -8106 244938
rect -8726 208938 -8694 209494
rect -8138 208938 -8106 209494
rect -8726 173494 -8106 208938
rect -8726 172938 -8694 173494
rect -8138 172938 -8106 173494
rect -8726 137494 -8106 172938
rect -8726 136938 -8694 137494
rect -8138 136938 -8106 137494
rect -8726 101494 -8106 136938
rect -8726 100938 -8694 101494
rect -8138 100938 -8106 101494
rect -8726 65494 -8106 100938
rect -8726 64938 -8694 65494
rect -8138 64938 -8106 65494
rect -8726 29494 -8106 64938
rect -8726 28938 -8694 29494
rect -8138 28938 -8106 29494
rect -8726 -7066 -8106 28938
rect -7766 710598 -7146 710630
rect -7766 710042 -7734 710598
rect -7178 710042 -7146 710598
rect -7766 673774 -7146 710042
rect -7766 673218 -7734 673774
rect -7178 673218 -7146 673774
rect -7766 637774 -7146 673218
rect -7766 637218 -7734 637774
rect -7178 637218 -7146 637774
rect -7766 601774 -7146 637218
rect -7766 601218 -7734 601774
rect -7178 601218 -7146 601774
rect -7766 565774 -7146 601218
rect -7766 565218 -7734 565774
rect -7178 565218 -7146 565774
rect -7766 529774 -7146 565218
rect -7766 529218 -7734 529774
rect -7178 529218 -7146 529774
rect -7766 493774 -7146 529218
rect -7766 493218 -7734 493774
rect -7178 493218 -7146 493774
rect -7766 457774 -7146 493218
rect -7766 457218 -7734 457774
rect -7178 457218 -7146 457774
rect -7766 421774 -7146 457218
rect -7766 421218 -7734 421774
rect -7178 421218 -7146 421774
rect -7766 385774 -7146 421218
rect -7766 385218 -7734 385774
rect -7178 385218 -7146 385774
rect -7766 349774 -7146 385218
rect -7766 349218 -7734 349774
rect -7178 349218 -7146 349774
rect -7766 313774 -7146 349218
rect -7766 313218 -7734 313774
rect -7178 313218 -7146 313774
rect -7766 277774 -7146 313218
rect -7766 277218 -7734 277774
rect -7178 277218 -7146 277774
rect -7766 241774 -7146 277218
rect -7766 241218 -7734 241774
rect -7178 241218 -7146 241774
rect -7766 205774 -7146 241218
rect -7766 205218 -7734 205774
rect -7178 205218 -7146 205774
rect -7766 169774 -7146 205218
rect -7766 169218 -7734 169774
rect -7178 169218 -7146 169774
rect -7766 133774 -7146 169218
rect -7766 133218 -7734 133774
rect -7178 133218 -7146 133774
rect -7766 97774 -7146 133218
rect -7766 97218 -7734 97774
rect -7178 97218 -7146 97774
rect -7766 61774 -7146 97218
rect -7766 61218 -7734 61774
rect -7178 61218 -7146 61774
rect -7766 25774 -7146 61218
rect -7766 25218 -7734 25774
rect -7178 25218 -7146 25774
rect -7766 -6106 -7146 25218
rect -6806 709638 -6186 709670
rect -6806 709082 -6774 709638
rect -6218 709082 -6186 709638
rect -6806 670054 -6186 709082
rect -6806 669498 -6774 670054
rect -6218 669498 -6186 670054
rect -6806 634054 -6186 669498
rect -6806 633498 -6774 634054
rect -6218 633498 -6186 634054
rect -6806 598054 -6186 633498
rect -6806 597498 -6774 598054
rect -6218 597498 -6186 598054
rect -6806 562054 -6186 597498
rect -6806 561498 -6774 562054
rect -6218 561498 -6186 562054
rect -6806 526054 -6186 561498
rect -6806 525498 -6774 526054
rect -6218 525498 -6186 526054
rect -6806 490054 -6186 525498
rect -6806 489498 -6774 490054
rect -6218 489498 -6186 490054
rect -6806 454054 -6186 489498
rect -6806 453498 -6774 454054
rect -6218 453498 -6186 454054
rect -6806 418054 -6186 453498
rect -6806 417498 -6774 418054
rect -6218 417498 -6186 418054
rect -6806 382054 -6186 417498
rect -6806 381498 -6774 382054
rect -6218 381498 -6186 382054
rect -6806 346054 -6186 381498
rect -6806 345498 -6774 346054
rect -6218 345498 -6186 346054
rect -6806 310054 -6186 345498
rect -6806 309498 -6774 310054
rect -6218 309498 -6186 310054
rect -6806 274054 -6186 309498
rect -6806 273498 -6774 274054
rect -6218 273498 -6186 274054
rect -6806 238054 -6186 273498
rect -6806 237498 -6774 238054
rect -6218 237498 -6186 238054
rect -6806 202054 -6186 237498
rect -6806 201498 -6774 202054
rect -6218 201498 -6186 202054
rect -6806 166054 -6186 201498
rect -6806 165498 -6774 166054
rect -6218 165498 -6186 166054
rect -6806 130054 -6186 165498
rect -6806 129498 -6774 130054
rect -6218 129498 -6186 130054
rect -6806 94054 -6186 129498
rect -6806 93498 -6774 94054
rect -6218 93498 -6186 94054
rect -6806 58054 -6186 93498
rect -6806 57498 -6774 58054
rect -6218 57498 -6186 58054
rect -6806 22054 -6186 57498
rect -6806 21498 -6774 22054
rect -6218 21498 -6186 22054
rect -6806 -5146 -6186 21498
rect -5846 708678 -5226 708710
rect -5846 708122 -5814 708678
rect -5258 708122 -5226 708678
rect -5846 666334 -5226 708122
rect -5846 665778 -5814 666334
rect -5258 665778 -5226 666334
rect -5846 630334 -5226 665778
rect -5846 629778 -5814 630334
rect -5258 629778 -5226 630334
rect -5846 594334 -5226 629778
rect -5846 593778 -5814 594334
rect -5258 593778 -5226 594334
rect -5846 558334 -5226 593778
rect -5846 557778 -5814 558334
rect -5258 557778 -5226 558334
rect -5846 522334 -5226 557778
rect -5846 521778 -5814 522334
rect -5258 521778 -5226 522334
rect -5846 486334 -5226 521778
rect -5846 485778 -5814 486334
rect -5258 485778 -5226 486334
rect -5846 450334 -5226 485778
rect -5846 449778 -5814 450334
rect -5258 449778 -5226 450334
rect -5846 414334 -5226 449778
rect -5846 413778 -5814 414334
rect -5258 413778 -5226 414334
rect -5846 378334 -5226 413778
rect -5846 377778 -5814 378334
rect -5258 377778 -5226 378334
rect -5846 342334 -5226 377778
rect -5846 341778 -5814 342334
rect -5258 341778 -5226 342334
rect -5846 306334 -5226 341778
rect -5846 305778 -5814 306334
rect -5258 305778 -5226 306334
rect -5846 270334 -5226 305778
rect -5846 269778 -5814 270334
rect -5258 269778 -5226 270334
rect -5846 234334 -5226 269778
rect -5846 233778 -5814 234334
rect -5258 233778 -5226 234334
rect -5846 198334 -5226 233778
rect -5846 197778 -5814 198334
rect -5258 197778 -5226 198334
rect -5846 162334 -5226 197778
rect -5846 161778 -5814 162334
rect -5258 161778 -5226 162334
rect -5846 126334 -5226 161778
rect -5846 125778 -5814 126334
rect -5258 125778 -5226 126334
rect -5846 90334 -5226 125778
rect -5846 89778 -5814 90334
rect -5258 89778 -5226 90334
rect -5846 54334 -5226 89778
rect -5846 53778 -5814 54334
rect -5258 53778 -5226 54334
rect -5846 18334 -5226 53778
rect -5846 17778 -5814 18334
rect -5258 17778 -5226 18334
rect -5846 -4186 -5226 17778
rect -4886 707718 -4266 707750
rect -4886 707162 -4854 707718
rect -4298 707162 -4266 707718
rect -4886 698614 -4266 707162
rect -4886 698058 -4854 698614
rect -4298 698058 -4266 698614
rect -4886 662614 -4266 698058
rect -4886 662058 -4854 662614
rect -4298 662058 -4266 662614
rect -4886 626614 -4266 662058
rect -4886 626058 -4854 626614
rect -4298 626058 -4266 626614
rect -4886 590614 -4266 626058
rect -4886 590058 -4854 590614
rect -4298 590058 -4266 590614
rect -4886 554614 -4266 590058
rect -4886 554058 -4854 554614
rect -4298 554058 -4266 554614
rect -4886 518614 -4266 554058
rect -4886 518058 -4854 518614
rect -4298 518058 -4266 518614
rect -4886 482614 -4266 518058
rect -4886 482058 -4854 482614
rect -4298 482058 -4266 482614
rect -4886 446614 -4266 482058
rect -4886 446058 -4854 446614
rect -4298 446058 -4266 446614
rect -4886 410614 -4266 446058
rect -4886 410058 -4854 410614
rect -4298 410058 -4266 410614
rect -4886 374614 -4266 410058
rect -4886 374058 -4854 374614
rect -4298 374058 -4266 374614
rect -4886 338614 -4266 374058
rect -4886 338058 -4854 338614
rect -4298 338058 -4266 338614
rect -4886 302614 -4266 338058
rect -4886 302058 -4854 302614
rect -4298 302058 -4266 302614
rect -4886 266614 -4266 302058
rect -4886 266058 -4854 266614
rect -4298 266058 -4266 266614
rect -4886 230614 -4266 266058
rect -4886 230058 -4854 230614
rect -4298 230058 -4266 230614
rect -4886 194614 -4266 230058
rect -4886 194058 -4854 194614
rect -4298 194058 -4266 194614
rect -4886 158614 -4266 194058
rect -4886 158058 -4854 158614
rect -4298 158058 -4266 158614
rect -4886 122614 -4266 158058
rect -4886 122058 -4854 122614
rect -4298 122058 -4266 122614
rect -4886 86614 -4266 122058
rect -4886 86058 -4854 86614
rect -4298 86058 -4266 86614
rect -4886 50614 -4266 86058
rect -4886 50058 -4854 50614
rect -4298 50058 -4266 50614
rect -4886 14614 -4266 50058
rect -4886 14058 -4854 14614
rect -4298 14058 -4266 14614
rect -4886 -3226 -4266 14058
rect -3926 706758 -3306 706790
rect -3926 706202 -3894 706758
rect -3338 706202 -3306 706758
rect -3926 694894 -3306 706202
rect -3926 694338 -3894 694894
rect -3338 694338 -3306 694894
rect -3926 658894 -3306 694338
rect -3926 658338 -3894 658894
rect -3338 658338 -3306 658894
rect -3926 622894 -3306 658338
rect -3926 622338 -3894 622894
rect -3338 622338 -3306 622894
rect -3926 586894 -3306 622338
rect -3926 586338 -3894 586894
rect -3338 586338 -3306 586894
rect -3926 550894 -3306 586338
rect -3926 550338 -3894 550894
rect -3338 550338 -3306 550894
rect -3926 514894 -3306 550338
rect -3926 514338 -3894 514894
rect -3338 514338 -3306 514894
rect -3926 478894 -3306 514338
rect -3926 478338 -3894 478894
rect -3338 478338 -3306 478894
rect -3926 442894 -3306 478338
rect -3926 442338 -3894 442894
rect -3338 442338 -3306 442894
rect -3926 406894 -3306 442338
rect -3926 406338 -3894 406894
rect -3338 406338 -3306 406894
rect -3926 370894 -3306 406338
rect -3926 370338 -3894 370894
rect -3338 370338 -3306 370894
rect -3926 334894 -3306 370338
rect -3926 334338 -3894 334894
rect -3338 334338 -3306 334894
rect -3926 298894 -3306 334338
rect -3926 298338 -3894 298894
rect -3338 298338 -3306 298894
rect -3926 262894 -3306 298338
rect -3926 262338 -3894 262894
rect -3338 262338 -3306 262894
rect -3926 226894 -3306 262338
rect -3926 226338 -3894 226894
rect -3338 226338 -3306 226894
rect -3926 190894 -3306 226338
rect -3926 190338 -3894 190894
rect -3338 190338 -3306 190894
rect -3926 154894 -3306 190338
rect -3926 154338 -3894 154894
rect -3338 154338 -3306 154894
rect -3926 118894 -3306 154338
rect -3926 118338 -3894 118894
rect -3338 118338 -3306 118894
rect -3926 82894 -3306 118338
rect -3926 82338 -3894 82894
rect -3338 82338 -3306 82894
rect -3926 46894 -3306 82338
rect -3926 46338 -3894 46894
rect -3338 46338 -3306 46894
rect -3926 10894 -3306 46338
rect -3926 10338 -3894 10894
rect -3338 10338 -3306 10894
rect -3926 -2266 -3306 10338
rect -2966 705798 -2346 705830
rect -2966 705242 -2934 705798
rect -2378 705242 -2346 705798
rect -2966 691174 -2346 705242
rect -2966 690618 -2934 691174
rect -2378 690618 -2346 691174
rect -2966 655174 -2346 690618
rect -2966 654618 -2934 655174
rect -2378 654618 -2346 655174
rect -2966 619174 -2346 654618
rect -2966 618618 -2934 619174
rect -2378 618618 -2346 619174
rect -2966 583174 -2346 618618
rect -2966 582618 -2934 583174
rect -2378 582618 -2346 583174
rect -2966 547174 -2346 582618
rect -2966 546618 -2934 547174
rect -2378 546618 -2346 547174
rect -2966 511174 -2346 546618
rect -2966 510618 -2934 511174
rect -2378 510618 -2346 511174
rect -2966 475174 -2346 510618
rect -2966 474618 -2934 475174
rect -2378 474618 -2346 475174
rect -2966 439174 -2346 474618
rect -2966 438618 -2934 439174
rect -2378 438618 -2346 439174
rect -2966 403174 -2346 438618
rect -2966 402618 -2934 403174
rect -2378 402618 -2346 403174
rect -2966 367174 -2346 402618
rect -2966 366618 -2934 367174
rect -2378 366618 -2346 367174
rect -2966 331174 -2346 366618
rect -2966 330618 -2934 331174
rect -2378 330618 -2346 331174
rect -2966 295174 -2346 330618
rect -2966 294618 -2934 295174
rect -2378 294618 -2346 295174
rect -2966 259174 -2346 294618
rect -2966 258618 -2934 259174
rect -2378 258618 -2346 259174
rect -2966 223174 -2346 258618
rect -2966 222618 -2934 223174
rect -2378 222618 -2346 223174
rect -2966 187174 -2346 222618
rect -2966 186618 -2934 187174
rect -2378 186618 -2346 187174
rect -2966 151174 -2346 186618
rect -2966 150618 -2934 151174
rect -2378 150618 -2346 151174
rect -2966 115174 -2346 150618
rect -2966 114618 -2934 115174
rect -2378 114618 -2346 115174
rect -2966 79174 -2346 114618
rect -2966 78618 -2934 79174
rect -2378 78618 -2346 79174
rect -2966 43174 -2346 78618
rect -2966 42618 -2934 43174
rect -2378 42618 -2346 43174
rect -2966 7174 -2346 42618
rect -2966 6618 -2934 7174
rect -2378 6618 -2346 7174
rect -2966 -1306 -2346 6618
rect -2006 704838 -1386 704870
rect -2006 704282 -1974 704838
rect -1418 704282 -1386 704838
rect -2006 687454 -1386 704282
rect -2006 686898 -1974 687454
rect -1418 686898 -1386 687454
rect -2006 651454 -1386 686898
rect -2006 650898 -1974 651454
rect -1418 650898 -1386 651454
rect -2006 615454 -1386 650898
rect -2006 614898 -1974 615454
rect -1418 614898 -1386 615454
rect -2006 579454 -1386 614898
rect -2006 578898 -1974 579454
rect -1418 578898 -1386 579454
rect -2006 543454 -1386 578898
rect -2006 542898 -1974 543454
rect -1418 542898 -1386 543454
rect -2006 507454 -1386 542898
rect -2006 506898 -1974 507454
rect -1418 506898 -1386 507454
rect -2006 471454 -1386 506898
rect -2006 470898 -1974 471454
rect -1418 470898 -1386 471454
rect -2006 435454 -1386 470898
rect -2006 434898 -1974 435454
rect -1418 434898 -1386 435454
rect -2006 399454 -1386 434898
rect -2006 398898 -1974 399454
rect -1418 398898 -1386 399454
rect -2006 363454 -1386 398898
rect -2006 362898 -1974 363454
rect -1418 362898 -1386 363454
rect -2006 327454 -1386 362898
rect -2006 326898 -1974 327454
rect -1418 326898 -1386 327454
rect -2006 291454 -1386 326898
rect -2006 290898 -1974 291454
rect -1418 290898 -1386 291454
rect -2006 255454 -1386 290898
rect -2006 254898 -1974 255454
rect -1418 254898 -1386 255454
rect -2006 219454 -1386 254898
rect -2006 218898 -1974 219454
rect -1418 218898 -1386 219454
rect -2006 183454 -1386 218898
rect -2006 182898 -1974 183454
rect -1418 182898 -1386 183454
rect -2006 147454 -1386 182898
rect -2006 146898 -1974 147454
rect -1418 146898 -1386 147454
rect -2006 111454 -1386 146898
rect -2006 110898 -1974 111454
rect -1418 110898 -1386 111454
rect -2006 75454 -1386 110898
rect -2006 74898 -1974 75454
rect -1418 74898 -1386 75454
rect -2006 39454 -1386 74898
rect -2006 38898 -1974 39454
rect -1418 38898 -1386 39454
rect -2006 3454 -1386 38898
rect -2006 2898 -1974 3454
rect -1418 2898 -1386 3454
rect -2006 -346 -1386 2898
rect -2006 -902 -1974 -346
rect -1418 -902 -1386 -346
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704282 1826 704838
rect 2382 704282 2414 704838
rect 1794 687454 2414 704282
rect 1794 686898 1826 687454
rect 2382 686898 2414 687454
rect 1794 651454 2414 686898
rect 1794 650898 1826 651454
rect 2382 650898 2414 651454
rect 1794 615454 2414 650898
rect 1794 614898 1826 615454
rect 2382 614898 2414 615454
rect 1794 579454 2414 614898
rect 1794 578898 1826 579454
rect 2382 578898 2414 579454
rect 1794 543454 2414 578898
rect 1794 542898 1826 543454
rect 2382 542898 2414 543454
rect 1794 507454 2414 542898
rect 1794 506898 1826 507454
rect 2382 506898 2414 507454
rect 1794 471454 2414 506898
rect 1794 470898 1826 471454
rect 2382 470898 2414 471454
rect 1794 435454 2414 470898
rect 1794 434898 1826 435454
rect 2382 434898 2414 435454
rect 1794 399454 2414 434898
rect 1794 398898 1826 399454
rect 2382 398898 2414 399454
rect 1794 363454 2414 398898
rect 1794 362898 1826 363454
rect 2382 362898 2414 363454
rect 1794 327454 2414 362898
rect 1794 326898 1826 327454
rect 2382 326898 2414 327454
rect 1794 291454 2414 326898
rect 1794 290898 1826 291454
rect 2382 290898 2414 291454
rect 1794 255454 2414 290898
rect 1794 254898 1826 255454
rect 2382 254898 2414 255454
rect 1794 219454 2414 254898
rect 1794 218898 1826 219454
rect 2382 218898 2414 219454
rect 1794 183454 2414 218898
rect 1794 182898 1826 183454
rect 2382 182898 2414 183454
rect 1794 147454 2414 182898
rect 1794 146898 1826 147454
rect 2382 146898 2414 147454
rect 1794 111454 2414 146898
rect 1794 110898 1826 111454
rect 2382 110898 2414 111454
rect 1794 75454 2414 110898
rect 1794 74898 1826 75454
rect 2382 74898 2414 75454
rect 1794 39454 2414 74898
rect 1794 38898 1826 39454
rect 2382 38898 2414 39454
rect 1794 3454 2414 38898
rect 1794 2898 1826 3454
rect 2382 2898 2414 3454
rect 1794 -346 2414 2898
rect 1794 -902 1826 -346
rect 2382 -902 2414 -346
rect -2966 -1862 -2934 -1306
rect -2378 -1862 -2346 -1306
rect -2966 -1894 -2346 -1862
rect -3926 -2822 -3894 -2266
rect -3338 -2822 -3306 -2266
rect -3926 -2854 -3306 -2822
rect -4886 -3782 -4854 -3226
rect -4298 -3782 -4266 -3226
rect -4886 -3814 -4266 -3782
rect -5846 -4742 -5814 -4186
rect -5258 -4742 -5226 -4186
rect -5846 -4774 -5226 -4742
rect -6806 -5702 -6774 -5146
rect -6218 -5702 -6186 -5146
rect -6806 -5734 -6186 -5702
rect -7766 -6662 -7734 -6106
rect -7178 -6662 -7146 -6106
rect -7766 -6694 -7146 -6662
rect -8726 -7622 -8694 -7066
rect -8138 -7622 -8106 -7066
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 5514 705798 6134 711590
rect 5514 705242 5546 705798
rect 6102 705242 6134 705798
rect 5514 691174 6134 705242
rect 5514 690618 5546 691174
rect 6102 690618 6134 691174
rect 5514 655174 6134 690618
rect 5514 654618 5546 655174
rect 6102 654618 6134 655174
rect 5514 619174 6134 654618
rect 5514 618618 5546 619174
rect 6102 618618 6134 619174
rect 5514 583174 6134 618618
rect 5514 582618 5546 583174
rect 6102 582618 6134 583174
rect 5514 547174 6134 582618
rect 5514 546618 5546 547174
rect 6102 546618 6134 547174
rect 5514 511174 6134 546618
rect 5514 510618 5546 511174
rect 6102 510618 6134 511174
rect 5514 475174 6134 510618
rect 5514 474618 5546 475174
rect 6102 474618 6134 475174
rect 5514 439174 6134 474618
rect 5514 438618 5546 439174
rect 6102 438618 6134 439174
rect 5514 403174 6134 438618
rect 5514 402618 5546 403174
rect 6102 402618 6134 403174
rect 5514 367174 6134 402618
rect 5514 366618 5546 367174
rect 6102 366618 6134 367174
rect 5514 331174 6134 366618
rect 5514 330618 5546 331174
rect 6102 330618 6134 331174
rect 5514 295174 6134 330618
rect 5514 294618 5546 295174
rect 6102 294618 6134 295174
rect 5514 259174 6134 294618
rect 5514 258618 5546 259174
rect 6102 258618 6134 259174
rect 5514 223174 6134 258618
rect 5514 222618 5546 223174
rect 6102 222618 6134 223174
rect 5514 187174 6134 222618
rect 5514 186618 5546 187174
rect 6102 186618 6134 187174
rect 5514 151174 6134 186618
rect 5514 150618 5546 151174
rect 6102 150618 6134 151174
rect 5514 115174 6134 150618
rect 5514 114618 5546 115174
rect 6102 114618 6134 115174
rect 5514 79174 6134 114618
rect 5514 78618 5546 79174
rect 6102 78618 6134 79174
rect 5514 43174 6134 78618
rect 5514 42618 5546 43174
rect 6102 42618 6134 43174
rect 5514 7174 6134 42618
rect 5514 6618 5546 7174
rect 6102 6618 6134 7174
rect 5514 -1306 6134 6618
rect 5514 -1862 5546 -1306
rect 6102 -1862 6134 -1306
rect 5514 -7654 6134 -1862
rect 9234 706758 9854 711590
rect 9234 706202 9266 706758
rect 9822 706202 9854 706758
rect 9234 694894 9854 706202
rect 9234 694338 9266 694894
rect 9822 694338 9854 694894
rect 9234 658894 9854 694338
rect 9234 658338 9266 658894
rect 9822 658338 9854 658894
rect 9234 622894 9854 658338
rect 9234 622338 9266 622894
rect 9822 622338 9854 622894
rect 9234 586894 9854 622338
rect 9234 586338 9266 586894
rect 9822 586338 9854 586894
rect 9234 550894 9854 586338
rect 9234 550338 9266 550894
rect 9822 550338 9854 550894
rect 9234 514894 9854 550338
rect 9234 514338 9266 514894
rect 9822 514338 9854 514894
rect 9234 478894 9854 514338
rect 9234 478338 9266 478894
rect 9822 478338 9854 478894
rect 9234 442894 9854 478338
rect 9234 442338 9266 442894
rect 9822 442338 9854 442894
rect 9234 406894 9854 442338
rect 9234 406338 9266 406894
rect 9822 406338 9854 406894
rect 9234 370894 9854 406338
rect 9234 370338 9266 370894
rect 9822 370338 9854 370894
rect 9234 334894 9854 370338
rect 9234 334338 9266 334894
rect 9822 334338 9854 334894
rect 9234 298894 9854 334338
rect 9234 298338 9266 298894
rect 9822 298338 9854 298894
rect 9234 262894 9854 298338
rect 9234 262338 9266 262894
rect 9822 262338 9854 262894
rect 9234 226894 9854 262338
rect 9234 226338 9266 226894
rect 9822 226338 9854 226894
rect 9234 190894 9854 226338
rect 9234 190338 9266 190894
rect 9822 190338 9854 190894
rect 9234 154894 9854 190338
rect 9234 154338 9266 154894
rect 9822 154338 9854 154894
rect 9234 118894 9854 154338
rect 9234 118338 9266 118894
rect 9822 118338 9854 118894
rect 9234 82894 9854 118338
rect 9234 82338 9266 82894
rect 9822 82338 9854 82894
rect 9234 46894 9854 82338
rect 9234 46338 9266 46894
rect 9822 46338 9854 46894
rect 9234 10894 9854 46338
rect 9234 10338 9266 10894
rect 9822 10338 9854 10894
rect 9234 -2266 9854 10338
rect 9234 -2822 9266 -2266
rect 9822 -2822 9854 -2266
rect 9234 -7654 9854 -2822
rect 12954 707718 13574 711590
rect 12954 707162 12986 707718
rect 13542 707162 13574 707718
rect 12954 698614 13574 707162
rect 12954 698058 12986 698614
rect 13542 698058 13574 698614
rect 12954 662614 13574 698058
rect 12954 662058 12986 662614
rect 13542 662058 13574 662614
rect 12954 626614 13574 662058
rect 12954 626058 12986 626614
rect 13542 626058 13574 626614
rect 12954 590614 13574 626058
rect 12954 590058 12986 590614
rect 13542 590058 13574 590614
rect 12954 554614 13574 590058
rect 12954 554058 12986 554614
rect 13542 554058 13574 554614
rect 12954 518614 13574 554058
rect 12954 518058 12986 518614
rect 13542 518058 13574 518614
rect 12954 482614 13574 518058
rect 12954 482058 12986 482614
rect 13542 482058 13574 482614
rect 12954 446614 13574 482058
rect 12954 446058 12986 446614
rect 13542 446058 13574 446614
rect 12954 410614 13574 446058
rect 12954 410058 12986 410614
rect 13542 410058 13574 410614
rect 12954 374614 13574 410058
rect 12954 374058 12986 374614
rect 13542 374058 13574 374614
rect 12954 338614 13574 374058
rect 12954 338058 12986 338614
rect 13542 338058 13574 338614
rect 12954 302614 13574 338058
rect 12954 302058 12986 302614
rect 13542 302058 13574 302614
rect 12954 266614 13574 302058
rect 12954 266058 12986 266614
rect 13542 266058 13574 266614
rect 12954 230614 13574 266058
rect 16674 708678 17294 711590
rect 16674 708122 16706 708678
rect 17262 708122 17294 708678
rect 16674 666334 17294 708122
rect 16674 665778 16706 666334
rect 17262 665778 17294 666334
rect 16674 630334 17294 665778
rect 16674 629778 16706 630334
rect 17262 629778 17294 630334
rect 16674 594334 17294 629778
rect 16674 593778 16706 594334
rect 17262 593778 17294 594334
rect 16674 558334 17294 593778
rect 16674 557778 16706 558334
rect 17262 557778 17294 558334
rect 16674 522334 17294 557778
rect 16674 521778 16706 522334
rect 17262 521778 17294 522334
rect 16674 486334 17294 521778
rect 16674 485778 16706 486334
rect 17262 485778 17294 486334
rect 16674 450334 17294 485778
rect 16674 449778 16706 450334
rect 17262 449778 17294 450334
rect 16674 414334 17294 449778
rect 16674 413778 16706 414334
rect 17262 413778 17294 414334
rect 16674 378334 17294 413778
rect 16674 377778 16706 378334
rect 17262 377778 17294 378334
rect 16674 342334 17294 377778
rect 16674 341778 16706 342334
rect 17262 341778 17294 342334
rect 16674 306334 17294 341778
rect 16674 305778 16706 306334
rect 17262 305778 17294 306334
rect 16674 270334 17294 305778
rect 16674 269778 16706 270334
rect 17262 269778 17294 270334
rect 16208 255454 16528 255486
rect 16208 255218 16250 255454
rect 16486 255218 16528 255454
rect 16208 255134 16528 255218
rect 16208 254898 16250 255134
rect 16486 254898 16528 255134
rect 16208 254866 16528 254898
rect 12954 230058 12986 230614
rect 13542 230058 13574 230614
rect 12954 194614 13574 230058
rect 16674 234334 17294 269778
rect 16674 233778 16706 234334
rect 17262 233778 17294 234334
rect 16208 219454 16528 219486
rect 16208 219218 16250 219454
rect 16486 219218 16528 219454
rect 16208 219134 16528 219218
rect 16208 218898 16250 219134
rect 16486 218898 16528 219134
rect 16208 218866 16528 218898
rect 12954 194058 12986 194614
rect 13542 194058 13574 194614
rect 12954 158614 13574 194058
rect 16674 198334 17294 233778
rect 16674 197778 16706 198334
rect 17262 197778 17294 198334
rect 16208 183454 16528 183486
rect 16208 183218 16250 183454
rect 16486 183218 16528 183454
rect 16208 183134 16528 183218
rect 16208 182898 16250 183134
rect 16486 182898 16528 183134
rect 16208 182866 16528 182898
rect 12954 158058 12986 158614
rect 13542 158058 13574 158614
rect 12954 122614 13574 158058
rect 16674 162334 17294 197778
rect 16674 161778 16706 162334
rect 17262 161778 17294 162334
rect 16674 149892 17294 161778
rect 20394 709638 21014 711590
rect 20394 709082 20426 709638
rect 20982 709082 21014 709638
rect 20394 670054 21014 709082
rect 20394 669498 20426 670054
rect 20982 669498 21014 670054
rect 20394 634054 21014 669498
rect 20394 633498 20426 634054
rect 20982 633498 21014 634054
rect 20394 598054 21014 633498
rect 20394 597498 20426 598054
rect 20982 597498 21014 598054
rect 20394 562054 21014 597498
rect 20394 561498 20426 562054
rect 20982 561498 21014 562054
rect 20394 526054 21014 561498
rect 20394 525498 20426 526054
rect 20982 525498 21014 526054
rect 20394 490054 21014 525498
rect 20394 489498 20426 490054
rect 20982 489498 21014 490054
rect 20394 454054 21014 489498
rect 20394 453498 20426 454054
rect 20982 453498 21014 454054
rect 20394 418054 21014 453498
rect 20394 417498 20426 418054
rect 20982 417498 21014 418054
rect 20394 382054 21014 417498
rect 20394 381498 20426 382054
rect 20982 381498 21014 382054
rect 20394 346054 21014 381498
rect 20394 345498 20426 346054
rect 20982 345498 21014 346054
rect 20394 310054 21014 345498
rect 20394 309498 20426 310054
rect 20982 309498 21014 310054
rect 20394 274054 21014 309498
rect 24114 710598 24734 711590
rect 24114 710042 24146 710598
rect 24702 710042 24734 710598
rect 24114 673774 24734 710042
rect 24114 673218 24146 673774
rect 24702 673218 24734 673774
rect 24114 637774 24734 673218
rect 24114 637218 24146 637774
rect 24702 637218 24734 637774
rect 24114 601774 24734 637218
rect 24114 601218 24146 601774
rect 24702 601218 24734 601774
rect 24114 565774 24734 601218
rect 24114 565218 24146 565774
rect 24702 565218 24734 565774
rect 24114 529774 24734 565218
rect 24114 529218 24146 529774
rect 24702 529218 24734 529774
rect 24114 493774 24734 529218
rect 24114 493218 24146 493774
rect 24702 493218 24734 493774
rect 24114 457774 24734 493218
rect 24114 457218 24146 457774
rect 24702 457218 24734 457774
rect 24114 421774 24734 457218
rect 24114 421218 24146 421774
rect 24702 421218 24734 421774
rect 24114 385774 24734 421218
rect 24114 385218 24146 385774
rect 24702 385218 24734 385774
rect 24114 349774 24734 385218
rect 24114 349218 24146 349774
rect 24702 349218 24734 349774
rect 24114 313774 24734 349218
rect 24114 313218 24146 313774
rect 24702 313218 24734 313774
rect 24114 282628 24734 313218
rect 27834 711558 28454 711590
rect 27834 711002 27866 711558
rect 28422 711002 28454 711558
rect 27834 677494 28454 711002
rect 27834 676938 27866 677494
rect 28422 676938 28454 677494
rect 27834 641494 28454 676938
rect 27834 640938 27866 641494
rect 28422 640938 28454 641494
rect 27834 605494 28454 640938
rect 27834 604938 27866 605494
rect 28422 604938 28454 605494
rect 27834 569494 28454 604938
rect 27834 568938 27866 569494
rect 28422 568938 28454 569494
rect 27834 533494 28454 568938
rect 27834 532938 27866 533494
rect 28422 532938 28454 533494
rect 27834 497494 28454 532938
rect 27834 496938 27866 497494
rect 28422 496938 28454 497494
rect 27834 461494 28454 496938
rect 27834 460938 27866 461494
rect 28422 460938 28454 461494
rect 27834 425494 28454 460938
rect 27834 424938 27866 425494
rect 28422 424938 28454 425494
rect 27834 389494 28454 424938
rect 27834 388938 27866 389494
rect 28422 388938 28454 389494
rect 27834 353494 28454 388938
rect 27834 352938 27866 353494
rect 28422 352938 28454 353494
rect 27834 317494 28454 352938
rect 27834 316938 27866 317494
rect 28422 316938 28454 317494
rect 20394 273498 20426 274054
rect 20982 273498 21014 274054
rect 20394 238054 21014 273498
rect 27834 281494 28454 316938
rect 27834 280938 27866 281494
rect 28422 280938 28454 281494
rect 23888 259174 24208 259206
rect 23888 258938 23930 259174
rect 24166 258938 24208 259174
rect 23888 258854 24208 258938
rect 23888 258618 23930 258854
rect 24166 258618 24208 258854
rect 23888 258586 24208 258618
rect 20394 237498 20426 238054
rect 20982 237498 21014 238054
rect 20394 202054 21014 237498
rect 27834 245494 28454 280938
rect 37794 704838 38414 711590
rect 37794 704282 37826 704838
rect 38382 704282 38414 704838
rect 37794 687454 38414 704282
rect 37794 686898 37826 687454
rect 38382 686898 38414 687454
rect 37794 651454 38414 686898
rect 37794 650898 37826 651454
rect 38382 650898 38414 651454
rect 37794 615454 38414 650898
rect 37794 614898 37826 615454
rect 38382 614898 38414 615454
rect 37794 579454 38414 614898
rect 37794 578898 37826 579454
rect 38382 578898 38414 579454
rect 37794 543454 38414 578898
rect 37794 542898 37826 543454
rect 38382 542898 38414 543454
rect 37794 507454 38414 542898
rect 37794 506898 37826 507454
rect 38382 506898 38414 507454
rect 37794 471454 38414 506898
rect 37794 470898 37826 471454
rect 38382 470898 38414 471454
rect 37794 435454 38414 470898
rect 37794 434898 37826 435454
rect 38382 434898 38414 435454
rect 37794 399454 38414 434898
rect 37794 398898 37826 399454
rect 38382 398898 38414 399454
rect 37794 363454 38414 398898
rect 37794 362898 37826 363454
rect 38382 362898 38414 363454
rect 37794 327454 38414 362898
rect 37794 326898 37826 327454
rect 38382 326898 38414 327454
rect 37794 291454 38414 326898
rect 37794 290898 37826 291454
rect 38382 290898 38414 291454
rect 31568 270334 31888 270366
rect 31568 270098 31610 270334
rect 31846 270098 31888 270334
rect 31568 270014 31888 270098
rect 31568 269778 31610 270014
rect 31846 269778 31888 270014
rect 31568 269746 31888 269778
rect 27834 244938 27866 245494
rect 28422 244938 28454 245494
rect 23888 223174 24208 223206
rect 23888 222938 23930 223174
rect 24166 222938 24208 223174
rect 23888 222854 24208 222938
rect 23888 222618 23930 222854
rect 24166 222618 24208 222854
rect 23888 222586 24208 222618
rect 20394 201498 20426 202054
rect 20982 201498 21014 202054
rect 20394 166054 21014 201498
rect 27834 209494 28454 244938
rect 37794 255454 38414 290898
rect 41514 705798 42134 711590
rect 41514 705242 41546 705798
rect 42102 705242 42134 705798
rect 41514 691174 42134 705242
rect 41514 690618 41546 691174
rect 42102 690618 42134 691174
rect 41514 655174 42134 690618
rect 41514 654618 41546 655174
rect 42102 654618 42134 655174
rect 41514 619174 42134 654618
rect 41514 618618 41546 619174
rect 42102 618618 42134 619174
rect 41514 583174 42134 618618
rect 41514 582618 41546 583174
rect 42102 582618 42134 583174
rect 41514 547174 42134 582618
rect 41514 546618 41546 547174
rect 42102 546618 42134 547174
rect 41514 511174 42134 546618
rect 41514 510618 41546 511174
rect 42102 510618 42134 511174
rect 41514 475174 42134 510618
rect 41514 474618 41546 475174
rect 42102 474618 42134 475174
rect 41514 439174 42134 474618
rect 41514 438618 41546 439174
rect 42102 438618 42134 439174
rect 41514 403174 42134 438618
rect 41514 402618 41546 403174
rect 42102 402618 42134 403174
rect 41514 367174 42134 402618
rect 41514 366618 41546 367174
rect 42102 366618 42134 367174
rect 41514 331174 42134 366618
rect 41514 330618 41546 331174
rect 42102 330618 42134 331174
rect 41514 295174 42134 330618
rect 41514 294618 41546 295174
rect 42102 294618 42134 295174
rect 39248 274054 39568 274086
rect 39248 273818 39290 274054
rect 39526 273818 39568 274054
rect 39248 273734 39568 273818
rect 39248 273498 39290 273734
rect 39526 273498 39568 273734
rect 39248 273466 39568 273498
rect 37794 254898 37826 255454
rect 38382 254898 38414 255454
rect 31568 234334 31888 234366
rect 31568 234098 31610 234334
rect 31846 234098 31888 234334
rect 31568 234014 31888 234098
rect 31568 233778 31610 234014
rect 31846 233778 31888 234014
rect 31568 233746 31888 233778
rect 27834 208938 27866 209494
rect 28422 208938 28454 209494
rect 23888 187174 24208 187206
rect 23888 186938 23930 187174
rect 24166 186938 24208 187174
rect 23888 186854 24208 186938
rect 23888 186618 23930 186854
rect 24166 186618 24208 186854
rect 23888 186586 24208 186618
rect 20394 165498 20426 166054
rect 20982 165498 21014 166054
rect 16208 147454 16528 147486
rect 16208 147218 16250 147454
rect 16486 147218 16528 147454
rect 16208 147134 16528 147218
rect 16208 146898 16250 147134
rect 16486 146898 16528 147134
rect 16208 146866 16528 146898
rect 12954 122058 12986 122614
rect 13542 122058 13574 122614
rect 12954 86614 13574 122058
rect 20394 130054 21014 165498
rect 27834 173494 28454 208938
rect 37794 219454 38414 254898
rect 41514 259174 42134 294618
rect 41514 258618 41546 259174
rect 42102 258618 42134 259174
rect 39248 238054 39568 238086
rect 39248 237818 39290 238054
rect 39526 237818 39568 238054
rect 39248 237734 39568 237818
rect 39248 237498 39290 237734
rect 39526 237498 39568 237734
rect 39248 237466 39568 237498
rect 37794 218898 37826 219454
rect 38382 218898 38414 219454
rect 31568 198334 31888 198366
rect 31568 198098 31610 198334
rect 31846 198098 31888 198334
rect 31568 198014 31888 198098
rect 31568 197778 31610 198014
rect 31846 197778 31888 198014
rect 31568 197746 31888 197778
rect 27834 172938 27866 173494
rect 28422 172938 28454 173494
rect 23888 151174 24208 151206
rect 23888 150938 23930 151174
rect 24166 150938 24208 151174
rect 23888 150854 24208 150938
rect 23888 150618 23930 150854
rect 24166 150618 24208 150854
rect 23888 150586 24208 150618
rect 20394 129498 20426 130054
rect 20982 129498 21014 130054
rect 17268 115174 17588 115206
rect 17268 114938 17310 115174
rect 17546 114938 17588 115174
rect 17268 114854 17588 114938
rect 17268 114618 17310 114854
rect 17546 114618 17588 114854
rect 17268 114586 17588 114618
rect 16208 111454 16528 111486
rect 16208 111218 16250 111454
rect 16486 111218 16528 111454
rect 16208 111134 16528 111218
rect 16208 110898 16250 111134
rect 16486 110898 16528 111134
rect 16208 110866 16528 110898
rect 12954 86058 12986 86614
rect 13542 86058 13574 86614
rect 12954 50614 13574 86058
rect 20394 94054 21014 129498
rect 27834 137494 28454 172938
rect 37794 183454 38414 218898
rect 41514 223174 42134 258618
rect 41514 222618 41546 223174
rect 42102 222618 42134 223174
rect 39248 202054 39568 202086
rect 39248 201818 39290 202054
rect 39526 201818 39568 202054
rect 39248 201734 39568 201818
rect 39248 201498 39290 201734
rect 39526 201498 39568 201734
rect 39248 201466 39568 201498
rect 37794 182898 37826 183454
rect 38382 182898 38414 183454
rect 31568 162334 31888 162366
rect 31568 162098 31610 162334
rect 31846 162098 31888 162334
rect 31568 162014 31888 162098
rect 31568 161778 31610 162014
rect 31846 161778 31888 162014
rect 31568 161746 31888 161778
rect 27834 136938 27866 137494
rect 28422 136938 28454 137494
rect 23888 115174 24208 115206
rect 23888 114938 23930 115174
rect 24166 114938 24208 115174
rect 23888 114854 24208 114938
rect 23888 114618 23930 114854
rect 24166 114618 24208 114854
rect 23888 114586 24208 114618
rect 20394 93498 20426 94054
rect 20982 93498 21014 94054
rect 17268 79174 17588 79206
rect 17268 78938 17310 79174
rect 17546 78938 17588 79174
rect 17268 78854 17588 78938
rect 17268 78618 17310 78854
rect 17546 78618 17588 78854
rect 17268 78586 17588 78618
rect 16208 75454 16528 75486
rect 16208 75218 16250 75454
rect 16486 75218 16528 75454
rect 16208 75134 16528 75218
rect 16208 74898 16250 75134
rect 16486 74898 16528 75134
rect 16208 74866 16528 74898
rect 12954 50058 12986 50614
rect 13542 50058 13574 50614
rect 12954 14614 13574 50058
rect 20394 58054 21014 93498
rect 27834 101494 28454 136938
rect 37794 147454 38414 182898
rect 41514 187174 42134 222618
rect 41514 186618 41546 187174
rect 42102 186618 42134 187174
rect 39248 166054 39568 166086
rect 39248 165818 39290 166054
rect 39526 165818 39568 166054
rect 39248 165734 39568 165818
rect 39248 165498 39290 165734
rect 39526 165498 39568 165734
rect 39248 165466 39568 165498
rect 37794 146898 37826 147454
rect 38382 146898 38414 147454
rect 31568 126334 31888 126366
rect 31568 126098 31610 126334
rect 31846 126098 31888 126334
rect 31568 126014 31888 126098
rect 31568 125778 31610 126014
rect 31846 125778 31888 126014
rect 31568 125746 31888 125778
rect 27834 100938 27866 101494
rect 28422 100938 28454 101494
rect 23888 79174 24208 79206
rect 23888 78938 23930 79174
rect 24166 78938 24208 79174
rect 23888 78854 24208 78938
rect 23888 78618 23930 78854
rect 24166 78618 24208 78854
rect 23888 78586 24208 78618
rect 20394 57498 20426 58054
rect 20982 57498 21014 58054
rect 17268 43174 17588 43206
rect 17268 42938 17310 43174
rect 17546 42938 17588 43174
rect 17268 42854 17588 42938
rect 17268 42618 17310 42854
rect 17546 42618 17588 42854
rect 17268 42586 17588 42618
rect 16208 39454 16528 39486
rect 16208 39218 16250 39454
rect 16486 39218 16528 39454
rect 16208 39134 16528 39218
rect 16208 38898 16250 39134
rect 16486 38898 16528 39134
rect 16208 38866 16528 38898
rect 12954 14058 12986 14614
rect 13542 14058 13574 14614
rect 12954 -3226 13574 14058
rect 20394 22054 21014 57498
rect 27834 65494 28454 100938
rect 37794 111454 38414 146898
rect 41514 151174 42134 186618
rect 41514 150618 41546 151174
rect 42102 150618 42134 151174
rect 39248 130054 39568 130086
rect 39248 129818 39290 130054
rect 39526 129818 39568 130054
rect 39248 129734 39568 129818
rect 39248 129498 39290 129734
rect 39526 129498 39568 129734
rect 39248 129466 39568 129498
rect 37794 110898 37826 111454
rect 38382 110898 38414 111454
rect 31568 90334 31888 90366
rect 31568 90098 31610 90334
rect 31846 90098 31888 90334
rect 31568 90014 31888 90098
rect 31568 89778 31610 90014
rect 31846 89778 31888 90014
rect 31568 89746 31888 89778
rect 27834 64938 27866 65494
rect 28422 64938 28454 65494
rect 23888 43174 24208 43206
rect 23888 42938 23930 43174
rect 24166 42938 24208 43174
rect 23888 42854 24208 42938
rect 23888 42618 23930 42854
rect 24166 42618 24208 42854
rect 23888 42586 24208 42618
rect 20394 21498 20426 22054
rect 20982 21498 21014 22054
rect 17268 7174 17588 7206
rect 17268 6938 17310 7174
rect 17546 6938 17588 7174
rect 17268 6854 17588 6938
rect 17268 6618 17310 6854
rect 17546 6618 17588 6854
rect 17268 6586 17588 6618
rect 12954 -3782 12986 -3226
rect 13542 -3782 13574 -3226
rect 12954 -7654 13574 -3782
rect 16674 -4186 17294 4076
rect 16674 -4742 16706 -4186
rect 17262 -4742 17294 -4186
rect 16674 -7654 17294 -4742
rect 20394 -5146 21014 21498
rect 27834 29494 28454 64938
rect 37794 75454 38414 110898
rect 41514 115174 42134 150618
rect 41514 114618 41546 115174
rect 42102 114618 42134 115174
rect 39248 94054 39568 94086
rect 39248 93818 39290 94054
rect 39526 93818 39568 94054
rect 39248 93734 39568 93818
rect 39248 93498 39290 93734
rect 39526 93498 39568 93734
rect 39248 93466 39568 93498
rect 37794 74898 37826 75454
rect 38382 74898 38414 75454
rect 31568 54334 31888 54366
rect 31568 54098 31610 54334
rect 31846 54098 31888 54334
rect 31568 54014 31888 54098
rect 31568 53778 31610 54014
rect 31846 53778 31888 54014
rect 31568 53746 31888 53778
rect 27834 28938 27866 29494
rect 28422 28938 28454 29494
rect 23888 7174 24208 7206
rect 23888 6938 23930 7174
rect 24166 6938 24208 7174
rect 23888 6854 24208 6938
rect 23888 6618 23930 6854
rect 24166 6618 24208 6854
rect 23888 6586 24208 6618
rect 20394 -5702 20426 -5146
rect 20982 -5702 21014 -5146
rect 20394 -7654 21014 -5702
rect 24114 -6106 24734 2988
rect 24114 -6662 24146 -6106
rect 24702 -6662 24734 -6106
rect 24114 -7654 24734 -6662
rect 27834 -7066 28454 28938
rect 37794 39454 38414 74898
rect 41514 79174 42134 114618
rect 41514 78618 41546 79174
rect 42102 78618 42134 79174
rect 39248 58054 39568 58086
rect 39248 57818 39290 58054
rect 39526 57818 39568 58054
rect 39248 57734 39568 57818
rect 39248 57498 39290 57734
rect 39526 57498 39568 57734
rect 39248 57466 39568 57498
rect 37794 38898 37826 39454
rect 38382 38898 38414 39454
rect 31568 18334 31888 18366
rect 31568 18098 31610 18334
rect 31846 18098 31888 18334
rect 31568 18014 31888 18098
rect 31568 17778 31610 18014
rect 31846 17778 31888 18014
rect 31568 17746 31888 17778
rect 27834 -7622 27866 -7066
rect 28422 -7622 28454 -7066
rect 27834 -7654 28454 -7622
rect 37794 3454 38414 38898
rect 41514 43174 42134 78618
rect 41514 42618 41546 43174
rect 42102 42618 42134 43174
rect 39248 22054 39568 22086
rect 39248 21818 39290 22054
rect 39526 21818 39568 22054
rect 39248 21734 39568 21818
rect 39248 21498 39290 21734
rect 39526 21498 39568 21734
rect 39248 21466 39568 21498
rect 37794 2898 37826 3454
rect 38382 2898 38414 3454
rect 37794 -346 38414 2898
rect 37794 -902 37826 -346
rect 38382 -902 38414 -346
rect 37794 -7654 38414 -902
rect 41514 7174 42134 42618
rect 41514 6618 41546 7174
rect 42102 6618 42134 7174
rect 41514 -1306 42134 6618
rect 41514 -1862 41546 -1306
rect 42102 -1862 42134 -1306
rect 41514 -7654 42134 -1862
rect 45234 706758 45854 711590
rect 45234 706202 45266 706758
rect 45822 706202 45854 706758
rect 45234 694894 45854 706202
rect 45234 694338 45266 694894
rect 45822 694338 45854 694894
rect 45234 658894 45854 694338
rect 45234 658338 45266 658894
rect 45822 658338 45854 658894
rect 45234 622894 45854 658338
rect 45234 622338 45266 622894
rect 45822 622338 45854 622894
rect 45234 586894 45854 622338
rect 45234 586338 45266 586894
rect 45822 586338 45854 586894
rect 45234 550894 45854 586338
rect 45234 550338 45266 550894
rect 45822 550338 45854 550894
rect 45234 514894 45854 550338
rect 45234 514338 45266 514894
rect 45822 514338 45854 514894
rect 45234 478894 45854 514338
rect 45234 478338 45266 478894
rect 45822 478338 45854 478894
rect 45234 442894 45854 478338
rect 45234 442338 45266 442894
rect 45822 442338 45854 442894
rect 45234 406894 45854 442338
rect 45234 406338 45266 406894
rect 45822 406338 45854 406894
rect 45234 370894 45854 406338
rect 45234 370338 45266 370894
rect 45822 370338 45854 370894
rect 45234 334894 45854 370338
rect 45234 334338 45266 334894
rect 45822 334338 45854 334894
rect 45234 298894 45854 334338
rect 45234 298338 45266 298894
rect 45822 298338 45854 298894
rect 45234 262894 45854 298338
rect 45234 262338 45266 262894
rect 45822 262338 45854 262894
rect 45234 226894 45854 262338
rect 48954 707718 49574 711590
rect 48954 707162 48986 707718
rect 49542 707162 49574 707718
rect 48954 698614 49574 707162
rect 48954 698058 48986 698614
rect 49542 698058 49574 698614
rect 48954 662614 49574 698058
rect 48954 662058 48986 662614
rect 49542 662058 49574 662614
rect 48954 626614 49574 662058
rect 48954 626058 48986 626614
rect 49542 626058 49574 626614
rect 48954 590614 49574 626058
rect 48954 590058 48986 590614
rect 49542 590058 49574 590614
rect 48954 554614 49574 590058
rect 48954 554058 48986 554614
rect 49542 554058 49574 554614
rect 48954 518614 49574 554058
rect 48954 518058 48986 518614
rect 49542 518058 49574 518614
rect 48954 482614 49574 518058
rect 48954 482058 48986 482614
rect 49542 482058 49574 482614
rect 48954 446614 49574 482058
rect 48954 446058 48986 446614
rect 49542 446058 49574 446614
rect 48954 410614 49574 446058
rect 48954 410058 48986 410614
rect 49542 410058 49574 410614
rect 48954 374614 49574 410058
rect 48954 374058 48986 374614
rect 49542 374058 49574 374614
rect 48954 338614 49574 374058
rect 48954 338058 48986 338614
rect 49542 338058 49574 338614
rect 48954 302614 49574 338058
rect 48954 302058 48986 302614
rect 49542 302058 49574 302614
rect 48954 266614 49574 302058
rect 48954 266058 48986 266614
rect 49542 266058 49574 266614
rect 46928 255454 47248 255486
rect 46928 255218 46970 255454
rect 47206 255218 47248 255454
rect 46928 255134 47248 255218
rect 46928 254898 46970 255134
rect 47206 254898 47248 255134
rect 46928 254866 47248 254898
rect 45234 226338 45266 226894
rect 45822 226338 45854 226894
rect 45234 190894 45854 226338
rect 48954 230614 49574 266058
rect 48954 230058 48986 230614
rect 49542 230058 49574 230614
rect 46928 219454 47248 219486
rect 46928 219218 46970 219454
rect 47206 219218 47248 219454
rect 46928 219134 47248 219218
rect 46928 218898 46970 219134
rect 47206 218898 47248 219134
rect 46928 218866 47248 218898
rect 45234 190338 45266 190894
rect 45822 190338 45854 190894
rect 45234 154894 45854 190338
rect 48954 194614 49574 230058
rect 48954 194058 48986 194614
rect 49542 194058 49574 194614
rect 46928 183454 47248 183486
rect 46928 183218 46970 183454
rect 47206 183218 47248 183454
rect 46928 183134 47248 183218
rect 46928 182898 46970 183134
rect 47206 182898 47248 183134
rect 46928 182866 47248 182898
rect 45234 154338 45266 154894
rect 45822 154338 45854 154894
rect 45234 118894 45854 154338
rect 48954 158614 49574 194058
rect 48954 158058 48986 158614
rect 49542 158058 49574 158614
rect 46928 147454 47248 147486
rect 46928 147218 46970 147454
rect 47206 147218 47248 147454
rect 46928 147134 47248 147218
rect 46928 146898 46970 147134
rect 47206 146898 47248 147134
rect 46928 146866 47248 146898
rect 45234 118338 45266 118894
rect 45822 118338 45854 118894
rect 45234 82894 45854 118338
rect 48954 122614 49574 158058
rect 48954 122058 48986 122614
rect 49542 122058 49574 122614
rect 46928 111454 47248 111486
rect 46928 111218 46970 111454
rect 47206 111218 47248 111454
rect 46928 111134 47248 111218
rect 46928 110898 46970 111134
rect 47206 110898 47248 111134
rect 46928 110866 47248 110898
rect 45234 82338 45266 82894
rect 45822 82338 45854 82894
rect 45234 46894 45854 82338
rect 48954 86614 49574 122058
rect 48954 86058 48986 86614
rect 49542 86058 49574 86614
rect 46928 75454 47248 75486
rect 46928 75218 46970 75454
rect 47206 75218 47248 75454
rect 46928 75134 47248 75218
rect 46928 74898 46970 75134
rect 47206 74898 47248 75134
rect 46928 74866 47248 74898
rect 45234 46338 45266 46894
rect 45822 46338 45854 46894
rect 45234 10894 45854 46338
rect 48954 50614 49574 86058
rect 48954 50058 48986 50614
rect 49542 50058 49574 50614
rect 46928 39454 47248 39486
rect 46928 39218 46970 39454
rect 47206 39218 47248 39454
rect 46928 39134 47248 39218
rect 46928 38898 46970 39134
rect 47206 38898 47248 39134
rect 46928 38866 47248 38898
rect 45234 10338 45266 10894
rect 45822 10338 45854 10894
rect 45234 -2266 45854 10338
rect 45234 -2822 45266 -2266
rect 45822 -2822 45854 -2266
rect 45234 -7654 45854 -2822
rect 48954 14614 49574 50058
rect 48954 14058 48986 14614
rect 49542 14058 49574 14614
rect 48954 -3226 49574 14058
rect 48954 -3782 48986 -3226
rect 49542 -3782 49574 -3226
rect 48954 -7654 49574 -3782
rect 52674 708678 53294 711590
rect 52674 708122 52706 708678
rect 53262 708122 53294 708678
rect 52674 666334 53294 708122
rect 52674 665778 52706 666334
rect 53262 665778 53294 666334
rect 52674 630334 53294 665778
rect 52674 629778 52706 630334
rect 53262 629778 53294 630334
rect 52674 594334 53294 629778
rect 52674 593778 52706 594334
rect 53262 593778 53294 594334
rect 52674 558334 53294 593778
rect 52674 557778 52706 558334
rect 53262 557778 53294 558334
rect 52674 522334 53294 557778
rect 52674 521778 52706 522334
rect 53262 521778 53294 522334
rect 52674 486334 53294 521778
rect 52674 485778 52706 486334
rect 53262 485778 53294 486334
rect 52674 450334 53294 485778
rect 52674 449778 52706 450334
rect 53262 449778 53294 450334
rect 52674 414334 53294 449778
rect 52674 413778 52706 414334
rect 53262 413778 53294 414334
rect 52674 378334 53294 413778
rect 52674 377778 52706 378334
rect 53262 377778 53294 378334
rect 52674 342334 53294 377778
rect 52674 341778 52706 342334
rect 53262 341778 53294 342334
rect 52674 306334 53294 341778
rect 52674 305778 52706 306334
rect 53262 305778 53294 306334
rect 52674 270334 53294 305778
rect 52674 269778 52706 270334
rect 53262 269778 53294 270334
rect 52674 234334 53294 269778
rect 56394 709638 57014 711590
rect 56394 709082 56426 709638
rect 56982 709082 57014 709638
rect 56394 670054 57014 709082
rect 56394 669498 56426 670054
rect 56982 669498 57014 670054
rect 56394 634054 57014 669498
rect 56394 633498 56426 634054
rect 56982 633498 57014 634054
rect 56394 598054 57014 633498
rect 56394 597498 56426 598054
rect 56982 597498 57014 598054
rect 56394 562054 57014 597498
rect 56394 561498 56426 562054
rect 56982 561498 57014 562054
rect 56394 526054 57014 561498
rect 56394 525498 56426 526054
rect 56982 525498 57014 526054
rect 56394 490054 57014 525498
rect 56394 489498 56426 490054
rect 56982 489498 57014 490054
rect 56394 454054 57014 489498
rect 56394 453498 56426 454054
rect 56982 453498 57014 454054
rect 56394 418054 57014 453498
rect 56394 417498 56426 418054
rect 56982 417498 57014 418054
rect 56394 382054 57014 417498
rect 56394 381498 56426 382054
rect 56982 381498 57014 382054
rect 56394 346054 57014 381498
rect 56394 345498 56426 346054
rect 56982 345498 57014 346054
rect 56394 310054 57014 345498
rect 56394 309498 56426 310054
rect 56982 309498 57014 310054
rect 56394 274054 57014 309498
rect 56394 273498 56426 274054
rect 56982 273498 57014 274054
rect 54608 259174 54928 259206
rect 54608 258938 54650 259174
rect 54886 258938 54928 259174
rect 54608 258854 54928 258938
rect 54608 258618 54650 258854
rect 54886 258618 54928 258854
rect 54608 258586 54928 258618
rect 52674 233778 52706 234334
rect 53262 233778 53294 234334
rect 52674 198334 53294 233778
rect 56394 238054 57014 273498
rect 56394 237498 56426 238054
rect 56982 237498 57014 238054
rect 54608 223174 54928 223206
rect 54608 222938 54650 223174
rect 54886 222938 54928 223174
rect 54608 222854 54928 222938
rect 54608 222618 54650 222854
rect 54886 222618 54928 222854
rect 54608 222586 54928 222618
rect 52674 197778 52706 198334
rect 53262 197778 53294 198334
rect 52674 162334 53294 197778
rect 56394 202054 57014 237498
rect 56394 201498 56426 202054
rect 56982 201498 57014 202054
rect 54608 187174 54928 187206
rect 54608 186938 54650 187174
rect 54886 186938 54928 187174
rect 54608 186854 54928 186938
rect 54608 186618 54650 186854
rect 54886 186618 54928 186854
rect 54608 186586 54928 186618
rect 52674 161778 52706 162334
rect 53262 161778 53294 162334
rect 52674 126334 53294 161778
rect 56394 166054 57014 201498
rect 56394 165498 56426 166054
rect 56982 165498 57014 166054
rect 54608 151174 54928 151206
rect 54608 150938 54650 151174
rect 54886 150938 54928 151174
rect 54608 150854 54928 150938
rect 54608 150618 54650 150854
rect 54886 150618 54928 150854
rect 54608 150586 54928 150618
rect 52674 125778 52706 126334
rect 53262 125778 53294 126334
rect 52674 90334 53294 125778
rect 56394 130054 57014 165498
rect 56394 129498 56426 130054
rect 56982 129498 57014 130054
rect 54608 115174 54928 115206
rect 54608 114938 54650 115174
rect 54886 114938 54928 115174
rect 54608 114854 54928 114938
rect 54608 114618 54650 114854
rect 54886 114618 54928 114854
rect 54608 114586 54928 114618
rect 52674 89778 52706 90334
rect 53262 89778 53294 90334
rect 52674 54334 53294 89778
rect 56394 94054 57014 129498
rect 56394 93498 56426 94054
rect 56982 93498 57014 94054
rect 54608 79174 54928 79206
rect 54608 78938 54650 79174
rect 54886 78938 54928 79174
rect 54608 78854 54928 78938
rect 54608 78618 54650 78854
rect 54886 78618 54928 78854
rect 54608 78586 54928 78618
rect 52674 53778 52706 54334
rect 53262 53778 53294 54334
rect 52674 18334 53294 53778
rect 56394 58054 57014 93498
rect 56394 57498 56426 58054
rect 56982 57498 57014 58054
rect 54608 43174 54928 43206
rect 54608 42938 54650 43174
rect 54886 42938 54928 43174
rect 54608 42854 54928 42938
rect 54608 42618 54650 42854
rect 54886 42618 54928 42854
rect 54608 42586 54928 42618
rect 52674 17778 52706 18334
rect 53262 17778 53294 18334
rect 52674 -4186 53294 17778
rect 56394 22054 57014 57498
rect 56394 21498 56426 22054
rect 56982 21498 57014 22054
rect 54608 7174 54928 7206
rect 54608 6938 54650 7174
rect 54886 6938 54928 7174
rect 54608 6854 54928 6938
rect 54608 6618 54650 6854
rect 54886 6618 54928 6854
rect 54608 6586 54928 6618
rect 52674 -4742 52706 -4186
rect 53262 -4742 53294 -4186
rect 52674 -7654 53294 -4742
rect 56394 -5146 57014 21498
rect 56394 -5702 56426 -5146
rect 56982 -5702 57014 -5146
rect 56394 -7654 57014 -5702
rect 60114 710598 60734 711590
rect 60114 710042 60146 710598
rect 60702 710042 60734 710598
rect 60114 673774 60734 710042
rect 60114 673218 60146 673774
rect 60702 673218 60734 673774
rect 60114 637774 60734 673218
rect 60114 637218 60146 637774
rect 60702 637218 60734 637774
rect 60114 601774 60734 637218
rect 60114 601218 60146 601774
rect 60702 601218 60734 601774
rect 60114 565774 60734 601218
rect 60114 565218 60146 565774
rect 60702 565218 60734 565774
rect 60114 529774 60734 565218
rect 60114 529218 60146 529774
rect 60702 529218 60734 529774
rect 60114 493774 60734 529218
rect 60114 493218 60146 493774
rect 60702 493218 60734 493774
rect 60114 457774 60734 493218
rect 60114 457218 60146 457774
rect 60702 457218 60734 457774
rect 60114 421774 60734 457218
rect 60114 421218 60146 421774
rect 60702 421218 60734 421774
rect 60114 385774 60734 421218
rect 60114 385218 60146 385774
rect 60702 385218 60734 385774
rect 60114 349774 60734 385218
rect 60114 349218 60146 349774
rect 60702 349218 60734 349774
rect 60114 313774 60734 349218
rect 60114 313218 60146 313774
rect 60702 313218 60734 313774
rect 60114 277774 60734 313218
rect 60114 277218 60146 277774
rect 60702 277218 60734 277774
rect 60114 241774 60734 277218
rect 63834 711558 64454 711590
rect 63834 711002 63866 711558
rect 64422 711002 64454 711558
rect 63834 677494 64454 711002
rect 63834 676938 63866 677494
rect 64422 676938 64454 677494
rect 63834 641494 64454 676938
rect 63834 640938 63866 641494
rect 64422 640938 64454 641494
rect 63834 605494 64454 640938
rect 63834 604938 63866 605494
rect 64422 604938 64454 605494
rect 63834 569494 64454 604938
rect 63834 568938 63866 569494
rect 64422 568938 64454 569494
rect 63834 533494 64454 568938
rect 63834 532938 63866 533494
rect 64422 532938 64454 533494
rect 63834 497494 64454 532938
rect 63834 496938 63866 497494
rect 64422 496938 64454 497494
rect 63834 461494 64454 496938
rect 63834 460938 63866 461494
rect 64422 460938 64454 461494
rect 63834 425494 64454 460938
rect 63834 424938 63866 425494
rect 64422 424938 64454 425494
rect 63834 389494 64454 424938
rect 63834 388938 63866 389494
rect 64422 388938 64454 389494
rect 63834 353494 64454 388938
rect 63834 352938 63866 353494
rect 64422 352938 64454 353494
rect 63834 317494 64454 352938
rect 63834 316938 63866 317494
rect 64422 316938 64454 317494
rect 63834 281494 64454 316938
rect 63834 280938 63866 281494
rect 64422 280938 64454 281494
rect 62288 270334 62608 270366
rect 62288 270098 62330 270334
rect 62566 270098 62608 270334
rect 62288 270014 62608 270098
rect 62288 269778 62330 270014
rect 62566 269778 62608 270014
rect 62288 269746 62608 269778
rect 60114 241218 60146 241774
rect 60702 241218 60734 241774
rect 60114 205774 60734 241218
rect 63834 245494 64454 280938
rect 73794 704838 74414 711590
rect 73794 704282 73826 704838
rect 74382 704282 74414 704838
rect 73794 687454 74414 704282
rect 73794 686898 73826 687454
rect 74382 686898 74414 687454
rect 73794 651454 74414 686898
rect 73794 650898 73826 651454
rect 74382 650898 74414 651454
rect 73794 615454 74414 650898
rect 73794 614898 73826 615454
rect 74382 614898 74414 615454
rect 73794 579454 74414 614898
rect 73794 578898 73826 579454
rect 74382 578898 74414 579454
rect 73794 543454 74414 578898
rect 73794 542898 73826 543454
rect 74382 542898 74414 543454
rect 73794 507454 74414 542898
rect 73794 506898 73826 507454
rect 74382 506898 74414 507454
rect 73794 471454 74414 506898
rect 73794 470898 73826 471454
rect 74382 470898 74414 471454
rect 73794 435454 74414 470898
rect 73794 434898 73826 435454
rect 74382 434898 74414 435454
rect 73794 399454 74414 434898
rect 73794 398898 73826 399454
rect 74382 398898 74414 399454
rect 73794 363454 74414 398898
rect 73794 362898 73826 363454
rect 74382 362898 74414 363454
rect 73794 327454 74414 362898
rect 73794 326898 73826 327454
rect 74382 326898 74414 327454
rect 73794 291454 74414 326898
rect 73794 290898 73826 291454
rect 74382 290898 74414 291454
rect 69968 274054 70288 274086
rect 69968 273818 70010 274054
rect 70246 273818 70288 274054
rect 69968 273734 70288 273818
rect 69968 273498 70010 273734
rect 70246 273498 70288 273734
rect 69968 273466 70288 273498
rect 63834 244938 63866 245494
rect 64422 244938 64454 245494
rect 62288 234334 62608 234366
rect 62288 234098 62330 234334
rect 62566 234098 62608 234334
rect 62288 234014 62608 234098
rect 62288 233778 62330 234014
rect 62566 233778 62608 234014
rect 62288 233746 62608 233778
rect 60114 205218 60146 205774
rect 60702 205218 60734 205774
rect 60114 169774 60734 205218
rect 63834 209494 64454 244938
rect 73794 255454 74414 290898
rect 77514 705798 78134 711590
rect 77514 705242 77546 705798
rect 78102 705242 78134 705798
rect 77514 691174 78134 705242
rect 77514 690618 77546 691174
rect 78102 690618 78134 691174
rect 77514 655174 78134 690618
rect 77514 654618 77546 655174
rect 78102 654618 78134 655174
rect 77514 619174 78134 654618
rect 77514 618618 77546 619174
rect 78102 618618 78134 619174
rect 77514 583174 78134 618618
rect 77514 582618 77546 583174
rect 78102 582618 78134 583174
rect 77514 547174 78134 582618
rect 77514 546618 77546 547174
rect 78102 546618 78134 547174
rect 77514 511174 78134 546618
rect 77514 510618 77546 511174
rect 78102 510618 78134 511174
rect 77514 475174 78134 510618
rect 77514 474618 77546 475174
rect 78102 474618 78134 475174
rect 77514 439174 78134 474618
rect 77514 438618 77546 439174
rect 78102 438618 78134 439174
rect 77514 403174 78134 438618
rect 77514 402618 77546 403174
rect 78102 402618 78134 403174
rect 77514 367174 78134 402618
rect 77514 366618 77546 367174
rect 78102 366618 78134 367174
rect 77514 331174 78134 366618
rect 77514 330618 77546 331174
rect 78102 330618 78134 331174
rect 77514 295174 78134 330618
rect 77514 294618 77546 295174
rect 78102 294618 78134 295174
rect 77514 282628 78134 294618
rect 81234 706758 81854 711590
rect 81234 706202 81266 706758
rect 81822 706202 81854 706758
rect 81234 694894 81854 706202
rect 81234 694338 81266 694894
rect 81822 694338 81854 694894
rect 81234 658894 81854 694338
rect 81234 658338 81266 658894
rect 81822 658338 81854 658894
rect 81234 622894 81854 658338
rect 81234 622338 81266 622894
rect 81822 622338 81854 622894
rect 81234 586894 81854 622338
rect 81234 586338 81266 586894
rect 81822 586338 81854 586894
rect 81234 550894 81854 586338
rect 81234 550338 81266 550894
rect 81822 550338 81854 550894
rect 81234 514894 81854 550338
rect 81234 514338 81266 514894
rect 81822 514338 81854 514894
rect 81234 478894 81854 514338
rect 81234 478338 81266 478894
rect 81822 478338 81854 478894
rect 81234 442894 81854 478338
rect 81234 442338 81266 442894
rect 81822 442338 81854 442894
rect 81234 406894 81854 442338
rect 81234 406338 81266 406894
rect 81822 406338 81854 406894
rect 81234 370894 81854 406338
rect 81234 370338 81266 370894
rect 81822 370338 81854 370894
rect 81234 334894 81854 370338
rect 81234 334338 81266 334894
rect 81822 334338 81854 334894
rect 81234 298894 81854 334338
rect 81234 298338 81266 298894
rect 81822 298338 81854 298894
rect 81234 262894 81854 298338
rect 84954 707718 85574 711590
rect 84954 707162 84986 707718
rect 85542 707162 85574 707718
rect 84954 698614 85574 707162
rect 84954 698058 84986 698614
rect 85542 698058 85574 698614
rect 84954 662614 85574 698058
rect 84954 662058 84986 662614
rect 85542 662058 85574 662614
rect 84954 626614 85574 662058
rect 84954 626058 84986 626614
rect 85542 626058 85574 626614
rect 84954 590614 85574 626058
rect 84954 590058 84986 590614
rect 85542 590058 85574 590614
rect 84954 554614 85574 590058
rect 84954 554058 84986 554614
rect 85542 554058 85574 554614
rect 84954 518614 85574 554058
rect 84954 518058 84986 518614
rect 85542 518058 85574 518614
rect 84954 482614 85574 518058
rect 84954 482058 84986 482614
rect 85542 482058 85574 482614
rect 84954 446614 85574 482058
rect 84954 446058 84986 446614
rect 85542 446058 85574 446614
rect 84954 410614 85574 446058
rect 84954 410058 84986 410614
rect 85542 410058 85574 410614
rect 84954 374614 85574 410058
rect 84954 374058 84986 374614
rect 85542 374058 85574 374614
rect 84954 338614 85574 374058
rect 84954 338058 84986 338614
rect 85542 338058 85574 338614
rect 84954 302614 85574 338058
rect 84954 302058 84986 302614
rect 85542 302058 85574 302614
rect 84954 282628 85574 302058
rect 88674 708678 89294 711590
rect 88674 708122 88706 708678
rect 89262 708122 89294 708678
rect 88674 666334 89294 708122
rect 88674 665778 88706 666334
rect 89262 665778 89294 666334
rect 88674 630334 89294 665778
rect 88674 629778 88706 630334
rect 89262 629778 89294 630334
rect 88674 594334 89294 629778
rect 88674 593778 88706 594334
rect 89262 593778 89294 594334
rect 88674 558334 89294 593778
rect 88674 557778 88706 558334
rect 89262 557778 89294 558334
rect 88674 522334 89294 557778
rect 88674 521778 88706 522334
rect 89262 521778 89294 522334
rect 88674 486334 89294 521778
rect 88674 485778 88706 486334
rect 89262 485778 89294 486334
rect 88674 450334 89294 485778
rect 88674 449778 88706 450334
rect 89262 449778 89294 450334
rect 88674 414334 89294 449778
rect 88674 413778 88706 414334
rect 89262 413778 89294 414334
rect 88674 378334 89294 413778
rect 88674 377778 88706 378334
rect 89262 377778 89294 378334
rect 88674 342334 89294 377778
rect 88674 341778 88706 342334
rect 89262 341778 89294 342334
rect 88674 306334 89294 341778
rect 88674 305778 88706 306334
rect 89262 305778 89294 306334
rect 81234 262338 81266 262894
rect 81822 262338 81854 262894
rect 73794 254898 73826 255454
rect 74382 254898 74414 255454
rect 69968 238054 70288 238086
rect 69968 237818 70010 238054
rect 70246 237818 70288 238054
rect 69968 237734 70288 237818
rect 69968 237498 70010 237734
rect 70246 237498 70288 237734
rect 69968 237466 70288 237498
rect 63834 208938 63866 209494
rect 64422 208938 64454 209494
rect 62288 198334 62608 198366
rect 62288 198098 62330 198334
rect 62566 198098 62608 198334
rect 62288 198014 62608 198098
rect 62288 197778 62330 198014
rect 62566 197778 62608 198014
rect 62288 197746 62608 197778
rect 60114 169218 60146 169774
rect 60702 169218 60734 169774
rect 60114 133774 60734 169218
rect 63834 173494 64454 208938
rect 73794 219454 74414 254898
rect 77648 255454 77968 255486
rect 77648 255218 77690 255454
rect 77926 255218 77968 255454
rect 77648 255134 77968 255218
rect 77648 254898 77690 255134
rect 77926 254898 77968 255134
rect 77648 254866 77968 254898
rect 81234 226894 81854 262338
rect 88674 270334 89294 305778
rect 92394 709638 93014 711590
rect 92394 709082 92426 709638
rect 92982 709082 93014 709638
rect 92394 670054 93014 709082
rect 92394 669498 92426 670054
rect 92982 669498 93014 670054
rect 92394 634054 93014 669498
rect 92394 633498 92426 634054
rect 92982 633498 93014 634054
rect 92394 598054 93014 633498
rect 92394 597498 92426 598054
rect 92982 597498 93014 598054
rect 92394 562054 93014 597498
rect 92394 561498 92426 562054
rect 92982 561498 93014 562054
rect 92394 526054 93014 561498
rect 92394 525498 92426 526054
rect 92982 525498 93014 526054
rect 92394 490054 93014 525498
rect 92394 489498 92426 490054
rect 92982 489498 93014 490054
rect 92394 454054 93014 489498
rect 92394 453498 92426 454054
rect 92982 453498 93014 454054
rect 92394 418054 93014 453498
rect 92394 417498 92426 418054
rect 92982 417498 93014 418054
rect 92394 382054 93014 417498
rect 92394 381498 92426 382054
rect 92982 381498 93014 382054
rect 92394 346054 93014 381498
rect 92394 345498 92426 346054
rect 92982 345498 93014 346054
rect 92394 310054 93014 345498
rect 92394 309498 92426 310054
rect 92982 309498 93014 310054
rect 92394 282628 93014 309498
rect 96114 710598 96734 711590
rect 96114 710042 96146 710598
rect 96702 710042 96734 710598
rect 96114 673774 96734 710042
rect 96114 673218 96146 673774
rect 96702 673218 96734 673774
rect 96114 637774 96734 673218
rect 96114 637218 96146 637774
rect 96702 637218 96734 637774
rect 96114 601774 96734 637218
rect 96114 601218 96146 601774
rect 96702 601218 96734 601774
rect 96114 565774 96734 601218
rect 96114 565218 96146 565774
rect 96702 565218 96734 565774
rect 96114 529774 96734 565218
rect 96114 529218 96146 529774
rect 96702 529218 96734 529774
rect 96114 493774 96734 529218
rect 96114 493218 96146 493774
rect 96702 493218 96734 493774
rect 96114 457774 96734 493218
rect 96114 457218 96146 457774
rect 96702 457218 96734 457774
rect 96114 421774 96734 457218
rect 96114 421218 96146 421774
rect 96702 421218 96734 421774
rect 96114 385774 96734 421218
rect 96114 385218 96146 385774
rect 96702 385218 96734 385774
rect 96114 349774 96734 385218
rect 96114 349218 96146 349774
rect 96702 349218 96734 349774
rect 96114 313774 96734 349218
rect 96114 313218 96146 313774
rect 96702 313218 96734 313774
rect 96114 277774 96734 313218
rect 96114 277218 96146 277774
rect 96702 277218 96734 277774
rect 88674 269778 88706 270334
rect 89262 269778 89294 270334
rect 85328 259174 85648 259206
rect 85328 258938 85370 259174
rect 85606 258938 85648 259174
rect 85328 258854 85648 258938
rect 85328 258618 85370 258854
rect 85606 258618 85648 258854
rect 85328 258586 85648 258618
rect 81234 226338 81266 226894
rect 81822 226338 81854 226894
rect 73794 218898 73826 219454
rect 74382 218898 74414 219454
rect 69968 202054 70288 202086
rect 69968 201818 70010 202054
rect 70246 201818 70288 202054
rect 69968 201734 70288 201818
rect 69968 201498 70010 201734
rect 70246 201498 70288 201734
rect 69968 201466 70288 201498
rect 63834 172938 63866 173494
rect 64422 172938 64454 173494
rect 62288 162334 62608 162366
rect 62288 162098 62330 162334
rect 62566 162098 62608 162334
rect 62288 162014 62608 162098
rect 62288 161778 62330 162014
rect 62566 161778 62608 162014
rect 62288 161746 62608 161778
rect 60114 133218 60146 133774
rect 60702 133218 60734 133774
rect 60114 97774 60734 133218
rect 63834 137494 64454 172938
rect 73794 183454 74414 218898
rect 77648 219454 77968 219486
rect 77648 219218 77690 219454
rect 77926 219218 77968 219454
rect 77648 219134 77968 219218
rect 77648 218898 77690 219134
rect 77926 218898 77968 219134
rect 77648 218866 77968 218898
rect 81234 190894 81854 226338
rect 88674 234334 89294 269778
rect 93008 270334 93328 270366
rect 93008 270098 93050 270334
rect 93286 270098 93328 270334
rect 93008 270014 93328 270098
rect 93008 269778 93050 270014
rect 93286 269778 93328 270014
rect 93008 269746 93328 269778
rect 96114 241774 96734 277218
rect 96114 241218 96146 241774
rect 96702 241218 96734 241774
rect 88674 233778 88706 234334
rect 89262 233778 89294 234334
rect 85328 223174 85648 223206
rect 85328 222938 85370 223174
rect 85606 222938 85648 223174
rect 85328 222854 85648 222938
rect 85328 222618 85370 222854
rect 85606 222618 85648 222854
rect 85328 222586 85648 222618
rect 81234 190338 81266 190894
rect 81822 190338 81854 190894
rect 73794 182898 73826 183454
rect 74382 182898 74414 183454
rect 69968 166054 70288 166086
rect 69968 165818 70010 166054
rect 70246 165818 70288 166054
rect 69968 165734 70288 165818
rect 69968 165498 70010 165734
rect 70246 165498 70288 165734
rect 69968 165466 70288 165498
rect 63834 136938 63866 137494
rect 64422 136938 64454 137494
rect 62288 126334 62608 126366
rect 62288 126098 62330 126334
rect 62566 126098 62608 126334
rect 62288 126014 62608 126098
rect 62288 125778 62330 126014
rect 62566 125778 62608 126014
rect 62288 125746 62608 125778
rect 60114 97218 60146 97774
rect 60702 97218 60734 97774
rect 60114 61774 60734 97218
rect 63834 101494 64454 136938
rect 73794 147454 74414 182898
rect 77648 183454 77968 183486
rect 77648 183218 77690 183454
rect 77926 183218 77968 183454
rect 77648 183134 77968 183218
rect 77648 182898 77690 183134
rect 77926 182898 77968 183134
rect 77648 182866 77968 182898
rect 81234 154894 81854 190338
rect 88674 198334 89294 233778
rect 93008 234334 93328 234366
rect 93008 234098 93050 234334
rect 93286 234098 93328 234334
rect 93008 234014 93328 234098
rect 93008 233778 93050 234014
rect 93286 233778 93328 234014
rect 93008 233746 93328 233778
rect 96114 205774 96734 241218
rect 96114 205218 96146 205774
rect 96702 205218 96734 205774
rect 88674 197778 88706 198334
rect 89262 197778 89294 198334
rect 85328 187174 85648 187206
rect 85328 186938 85370 187174
rect 85606 186938 85648 187174
rect 85328 186854 85648 186938
rect 85328 186618 85370 186854
rect 85606 186618 85648 186854
rect 85328 186586 85648 186618
rect 81234 154338 81266 154894
rect 81822 154338 81854 154894
rect 73794 146898 73826 147454
rect 74382 146898 74414 147454
rect 69968 130054 70288 130086
rect 69968 129818 70010 130054
rect 70246 129818 70288 130054
rect 69968 129734 70288 129818
rect 69968 129498 70010 129734
rect 70246 129498 70288 129734
rect 69968 129466 70288 129498
rect 63834 100938 63866 101494
rect 64422 100938 64454 101494
rect 62288 90334 62608 90366
rect 62288 90098 62330 90334
rect 62566 90098 62608 90334
rect 62288 90014 62608 90098
rect 62288 89778 62330 90014
rect 62566 89778 62608 90014
rect 62288 89746 62608 89778
rect 60114 61218 60146 61774
rect 60702 61218 60734 61774
rect 60114 25774 60734 61218
rect 63834 65494 64454 100938
rect 73794 111454 74414 146898
rect 77648 147454 77968 147486
rect 77648 147218 77690 147454
rect 77926 147218 77968 147454
rect 77648 147134 77968 147218
rect 77648 146898 77690 147134
rect 77926 146898 77968 147134
rect 77648 146866 77968 146898
rect 81234 118894 81854 154338
rect 88674 162334 89294 197778
rect 93008 198334 93328 198366
rect 93008 198098 93050 198334
rect 93286 198098 93328 198334
rect 93008 198014 93328 198098
rect 93008 197778 93050 198014
rect 93286 197778 93328 198014
rect 93008 197746 93328 197778
rect 96114 169774 96734 205218
rect 96114 169218 96146 169774
rect 96702 169218 96734 169774
rect 88674 161778 88706 162334
rect 89262 161778 89294 162334
rect 85328 151174 85648 151206
rect 85328 150938 85370 151174
rect 85606 150938 85648 151174
rect 85328 150854 85648 150938
rect 85328 150618 85370 150854
rect 85606 150618 85648 150854
rect 85328 150586 85648 150618
rect 81234 118338 81266 118894
rect 81822 118338 81854 118894
rect 73794 110898 73826 111454
rect 74382 110898 74414 111454
rect 69968 94054 70288 94086
rect 69968 93818 70010 94054
rect 70246 93818 70288 94054
rect 69968 93734 70288 93818
rect 69968 93498 70010 93734
rect 70246 93498 70288 93734
rect 69968 93466 70288 93498
rect 63834 64938 63866 65494
rect 64422 64938 64454 65494
rect 62288 54334 62608 54366
rect 62288 54098 62330 54334
rect 62566 54098 62608 54334
rect 62288 54014 62608 54098
rect 62288 53778 62330 54014
rect 62566 53778 62608 54014
rect 62288 53746 62608 53778
rect 60114 25218 60146 25774
rect 60702 25218 60734 25774
rect 60114 -6106 60734 25218
rect 63834 29494 64454 64938
rect 73794 75454 74414 110898
rect 77648 111454 77968 111486
rect 77648 111218 77690 111454
rect 77926 111218 77968 111454
rect 77648 111134 77968 111218
rect 77648 110898 77690 111134
rect 77926 110898 77968 111134
rect 77648 110866 77968 110898
rect 81234 82894 81854 118338
rect 88674 126334 89294 161778
rect 93008 162334 93328 162366
rect 93008 162098 93050 162334
rect 93286 162098 93328 162334
rect 93008 162014 93328 162098
rect 93008 161778 93050 162014
rect 93286 161778 93328 162014
rect 93008 161746 93328 161778
rect 96114 133774 96734 169218
rect 96114 133218 96146 133774
rect 96702 133218 96734 133774
rect 88674 125778 88706 126334
rect 89262 125778 89294 126334
rect 85328 115174 85648 115206
rect 85328 114938 85370 115174
rect 85606 114938 85648 115174
rect 85328 114854 85648 114938
rect 85328 114618 85370 114854
rect 85606 114618 85648 114854
rect 85328 114586 85648 114618
rect 81234 82338 81266 82894
rect 81822 82338 81854 82894
rect 73794 74898 73826 75454
rect 74382 74898 74414 75454
rect 69968 58054 70288 58086
rect 69968 57818 70010 58054
rect 70246 57818 70288 58054
rect 69968 57734 70288 57818
rect 69968 57498 70010 57734
rect 70246 57498 70288 57734
rect 69968 57466 70288 57498
rect 63834 28938 63866 29494
rect 64422 28938 64454 29494
rect 62288 18334 62608 18366
rect 62288 18098 62330 18334
rect 62566 18098 62608 18334
rect 62288 18014 62608 18098
rect 62288 17778 62330 18014
rect 62566 17778 62608 18014
rect 62288 17746 62608 17778
rect 60114 -6662 60146 -6106
rect 60702 -6662 60734 -6106
rect 60114 -7654 60734 -6662
rect 63834 -7066 64454 28938
rect 73794 39454 74414 74898
rect 77648 75454 77968 75486
rect 77648 75218 77690 75454
rect 77926 75218 77968 75454
rect 77648 75134 77968 75218
rect 77648 74898 77690 75134
rect 77926 74898 77968 75134
rect 77648 74866 77968 74898
rect 81234 46894 81854 82338
rect 88674 90334 89294 125778
rect 93008 126334 93328 126366
rect 93008 126098 93050 126334
rect 93286 126098 93328 126334
rect 93008 126014 93328 126098
rect 93008 125778 93050 126014
rect 93286 125778 93328 126014
rect 93008 125746 93328 125778
rect 96114 97774 96734 133218
rect 96114 97218 96146 97774
rect 96702 97218 96734 97774
rect 88674 89778 88706 90334
rect 89262 89778 89294 90334
rect 85328 79174 85648 79206
rect 85328 78938 85370 79174
rect 85606 78938 85648 79174
rect 85328 78854 85648 78938
rect 85328 78618 85370 78854
rect 85606 78618 85648 78854
rect 85328 78586 85648 78618
rect 81234 46338 81266 46894
rect 81822 46338 81854 46894
rect 73794 38898 73826 39454
rect 74382 38898 74414 39454
rect 69968 22054 70288 22086
rect 69968 21818 70010 22054
rect 70246 21818 70288 22054
rect 69968 21734 70288 21818
rect 69968 21498 70010 21734
rect 70246 21498 70288 21734
rect 69968 21466 70288 21498
rect 63834 -7622 63866 -7066
rect 64422 -7622 64454 -7066
rect 63834 -7654 64454 -7622
rect 73794 3454 74414 38898
rect 77648 39454 77968 39486
rect 77648 39218 77690 39454
rect 77926 39218 77968 39454
rect 77648 39134 77968 39218
rect 77648 38898 77690 39134
rect 77926 38898 77968 39134
rect 77648 38866 77968 38898
rect 73794 2898 73826 3454
rect 74382 2898 74414 3454
rect 81234 10894 81854 46338
rect 88674 54334 89294 89778
rect 93008 90334 93328 90366
rect 93008 90098 93050 90334
rect 93286 90098 93328 90334
rect 93008 90014 93328 90098
rect 93008 89778 93050 90014
rect 93286 89778 93328 90014
rect 93008 89746 93328 89778
rect 96114 61774 96734 97218
rect 96114 61218 96146 61774
rect 96702 61218 96734 61774
rect 88674 53778 88706 54334
rect 89262 53778 89294 54334
rect 85328 43174 85648 43206
rect 85328 42938 85370 43174
rect 85606 42938 85648 43174
rect 85328 42854 85648 42938
rect 85328 42618 85370 42854
rect 85606 42618 85648 42854
rect 85328 42586 85648 42618
rect 81234 10338 81266 10894
rect 81822 10338 81854 10894
rect 73794 -346 74414 2898
rect 73794 -902 73826 -346
rect 74382 -902 74414 -346
rect 73794 -7654 74414 -902
rect 77514 -1306 78134 2988
rect 77514 -1862 77546 -1306
rect 78102 -1862 78134 -1306
rect 77514 -7654 78134 -1862
rect 81234 -2266 81854 10338
rect 88674 18334 89294 53778
rect 93008 54334 93328 54366
rect 93008 54098 93050 54334
rect 93286 54098 93328 54334
rect 93008 54014 93328 54098
rect 93008 53778 93050 54014
rect 93286 53778 93328 54014
rect 93008 53746 93328 53778
rect 96114 25774 96734 61218
rect 96114 25218 96146 25774
rect 96702 25218 96734 25774
rect 88674 17778 88706 18334
rect 89262 17778 89294 18334
rect 85328 7174 85648 7206
rect 85328 6938 85370 7174
rect 85606 6938 85648 7174
rect 85328 6854 85648 6938
rect 85328 6618 85370 6854
rect 85606 6618 85648 6854
rect 85328 6586 85648 6618
rect 81234 -2822 81266 -2266
rect 81822 -2822 81854 -2266
rect 81234 -7654 81854 -2822
rect 84954 -3226 85574 2988
rect 84954 -3782 84986 -3226
rect 85542 -3782 85574 -3226
rect 84954 -7654 85574 -3782
rect 88674 -4186 89294 17778
rect 93008 18334 93328 18366
rect 93008 18098 93050 18334
rect 93286 18098 93328 18334
rect 93008 18014 93328 18098
rect 93008 17778 93050 18014
rect 93286 17778 93328 18014
rect 93008 17746 93328 17778
rect 88674 -4742 88706 -4186
rect 89262 -4742 89294 -4186
rect 88674 -7654 89294 -4742
rect 92394 -5146 93014 2988
rect 92394 -5702 92426 -5146
rect 92982 -5702 93014 -5146
rect 92394 -7654 93014 -5702
rect 96114 -6106 96734 25218
rect 96114 -6662 96146 -6106
rect 96702 -6662 96734 -6106
rect 96114 -7654 96734 -6662
rect 99834 711558 100454 711590
rect 99834 711002 99866 711558
rect 100422 711002 100454 711558
rect 99834 677494 100454 711002
rect 99834 676938 99866 677494
rect 100422 676938 100454 677494
rect 99834 641494 100454 676938
rect 99834 640938 99866 641494
rect 100422 640938 100454 641494
rect 99834 605494 100454 640938
rect 99834 604938 99866 605494
rect 100422 604938 100454 605494
rect 99834 569494 100454 604938
rect 99834 568938 99866 569494
rect 100422 568938 100454 569494
rect 99834 533494 100454 568938
rect 99834 532938 99866 533494
rect 100422 532938 100454 533494
rect 99834 497494 100454 532938
rect 99834 496938 99866 497494
rect 100422 496938 100454 497494
rect 99834 461494 100454 496938
rect 99834 460938 99866 461494
rect 100422 460938 100454 461494
rect 99834 425494 100454 460938
rect 99834 424938 99866 425494
rect 100422 424938 100454 425494
rect 99834 389494 100454 424938
rect 99834 388938 99866 389494
rect 100422 388938 100454 389494
rect 99834 353494 100454 388938
rect 99834 352938 99866 353494
rect 100422 352938 100454 353494
rect 99834 317494 100454 352938
rect 99834 316938 99866 317494
rect 100422 316938 100454 317494
rect 99834 281494 100454 316938
rect 99834 280938 99866 281494
rect 100422 280938 100454 281494
rect 99834 245494 100454 280938
rect 109794 704838 110414 711590
rect 109794 704282 109826 704838
rect 110382 704282 110414 704838
rect 109794 687454 110414 704282
rect 109794 686898 109826 687454
rect 110382 686898 110414 687454
rect 109794 651454 110414 686898
rect 109794 650898 109826 651454
rect 110382 650898 110414 651454
rect 109794 615454 110414 650898
rect 109794 614898 109826 615454
rect 110382 614898 110414 615454
rect 109794 579454 110414 614898
rect 109794 578898 109826 579454
rect 110382 578898 110414 579454
rect 109794 543454 110414 578898
rect 109794 542898 109826 543454
rect 110382 542898 110414 543454
rect 109794 507454 110414 542898
rect 109794 506898 109826 507454
rect 110382 506898 110414 507454
rect 109794 471454 110414 506898
rect 109794 470898 109826 471454
rect 110382 470898 110414 471454
rect 109794 435454 110414 470898
rect 109794 434898 109826 435454
rect 110382 434898 110414 435454
rect 109794 399454 110414 434898
rect 109794 398898 109826 399454
rect 110382 398898 110414 399454
rect 109794 363454 110414 398898
rect 109794 362898 109826 363454
rect 110382 362898 110414 363454
rect 109794 327454 110414 362898
rect 109794 326898 109826 327454
rect 110382 326898 110414 327454
rect 109794 291454 110414 326898
rect 109794 290898 109826 291454
rect 110382 290898 110414 291454
rect 100688 274054 101008 274086
rect 100688 273818 100730 274054
rect 100966 273818 101008 274054
rect 100688 273734 101008 273818
rect 100688 273498 100730 273734
rect 100966 273498 101008 273734
rect 100688 273466 101008 273498
rect 108368 255454 108688 255486
rect 108368 255218 108410 255454
rect 108646 255218 108688 255454
rect 108368 255134 108688 255218
rect 108368 254898 108410 255134
rect 108646 254898 108688 255134
rect 108368 254866 108688 254898
rect 109794 255454 110414 290898
rect 109794 254898 109826 255454
rect 110382 254898 110414 255454
rect 99834 244938 99866 245494
rect 100422 244938 100454 245494
rect 99834 209494 100454 244938
rect 100688 238054 101008 238086
rect 100688 237818 100730 238054
rect 100966 237818 101008 238054
rect 100688 237734 101008 237818
rect 100688 237498 100730 237734
rect 100966 237498 101008 237734
rect 100688 237466 101008 237498
rect 108368 219454 108688 219486
rect 108368 219218 108410 219454
rect 108646 219218 108688 219454
rect 108368 219134 108688 219218
rect 108368 218898 108410 219134
rect 108646 218898 108688 219134
rect 108368 218866 108688 218898
rect 109794 219454 110414 254898
rect 109794 218898 109826 219454
rect 110382 218898 110414 219454
rect 99834 208938 99866 209494
rect 100422 208938 100454 209494
rect 99834 173494 100454 208938
rect 100688 202054 101008 202086
rect 100688 201818 100730 202054
rect 100966 201818 101008 202054
rect 100688 201734 101008 201818
rect 100688 201498 100730 201734
rect 100966 201498 101008 201734
rect 100688 201466 101008 201498
rect 108368 183454 108688 183486
rect 108368 183218 108410 183454
rect 108646 183218 108688 183454
rect 108368 183134 108688 183218
rect 108368 182898 108410 183134
rect 108646 182898 108688 183134
rect 108368 182866 108688 182898
rect 109794 183454 110414 218898
rect 109794 182898 109826 183454
rect 110382 182898 110414 183454
rect 99834 172938 99866 173494
rect 100422 172938 100454 173494
rect 99834 137494 100454 172938
rect 100688 166054 101008 166086
rect 100688 165818 100730 166054
rect 100966 165818 101008 166054
rect 100688 165734 101008 165818
rect 100688 165498 100730 165734
rect 100966 165498 101008 165734
rect 100688 165466 101008 165498
rect 108368 147454 108688 147486
rect 108368 147218 108410 147454
rect 108646 147218 108688 147454
rect 108368 147134 108688 147218
rect 108368 146898 108410 147134
rect 108646 146898 108688 147134
rect 108368 146866 108688 146898
rect 109794 147454 110414 182898
rect 109794 146898 109826 147454
rect 110382 146898 110414 147454
rect 99834 136938 99866 137494
rect 100422 136938 100454 137494
rect 99834 101494 100454 136938
rect 100688 130054 101008 130086
rect 100688 129818 100730 130054
rect 100966 129818 101008 130054
rect 100688 129734 101008 129818
rect 100688 129498 100730 129734
rect 100966 129498 101008 129734
rect 100688 129466 101008 129498
rect 108368 111454 108688 111486
rect 108368 111218 108410 111454
rect 108646 111218 108688 111454
rect 108368 111134 108688 111218
rect 108368 110898 108410 111134
rect 108646 110898 108688 111134
rect 108368 110866 108688 110898
rect 109794 111454 110414 146898
rect 113514 705798 114134 711590
rect 113514 705242 113546 705798
rect 114102 705242 114134 705798
rect 113514 691174 114134 705242
rect 113514 690618 113546 691174
rect 114102 690618 114134 691174
rect 113514 655174 114134 690618
rect 113514 654618 113546 655174
rect 114102 654618 114134 655174
rect 113514 619174 114134 654618
rect 113514 618618 113546 619174
rect 114102 618618 114134 619174
rect 113514 583174 114134 618618
rect 113514 582618 113546 583174
rect 114102 582618 114134 583174
rect 113514 547174 114134 582618
rect 113514 546618 113546 547174
rect 114102 546618 114134 547174
rect 113514 511174 114134 546618
rect 113514 510618 113546 511174
rect 114102 510618 114134 511174
rect 113514 475174 114134 510618
rect 113514 474618 113546 475174
rect 114102 474618 114134 475174
rect 113514 439174 114134 474618
rect 113514 438618 113546 439174
rect 114102 438618 114134 439174
rect 113514 403174 114134 438618
rect 113514 402618 113546 403174
rect 114102 402618 114134 403174
rect 113514 367174 114134 402618
rect 113514 366618 113546 367174
rect 114102 366618 114134 367174
rect 113514 331174 114134 366618
rect 113514 330618 113546 331174
rect 114102 330618 114134 331174
rect 113514 295174 114134 330618
rect 113514 294618 113546 295174
rect 114102 294618 114134 295174
rect 113514 259174 114134 294618
rect 117234 706758 117854 711590
rect 117234 706202 117266 706758
rect 117822 706202 117854 706758
rect 117234 694894 117854 706202
rect 117234 694338 117266 694894
rect 117822 694338 117854 694894
rect 117234 658894 117854 694338
rect 117234 658338 117266 658894
rect 117822 658338 117854 658894
rect 117234 622894 117854 658338
rect 117234 622338 117266 622894
rect 117822 622338 117854 622894
rect 117234 586894 117854 622338
rect 117234 586338 117266 586894
rect 117822 586338 117854 586894
rect 117234 550894 117854 586338
rect 117234 550338 117266 550894
rect 117822 550338 117854 550894
rect 117234 514894 117854 550338
rect 117234 514338 117266 514894
rect 117822 514338 117854 514894
rect 117234 478894 117854 514338
rect 117234 478338 117266 478894
rect 117822 478338 117854 478894
rect 117234 442894 117854 478338
rect 117234 442338 117266 442894
rect 117822 442338 117854 442894
rect 117234 406894 117854 442338
rect 117234 406338 117266 406894
rect 117822 406338 117854 406894
rect 117234 370894 117854 406338
rect 117234 370338 117266 370894
rect 117822 370338 117854 370894
rect 117234 334894 117854 370338
rect 117234 334338 117266 334894
rect 117822 334338 117854 334894
rect 117234 298894 117854 334338
rect 117234 298338 117266 298894
rect 117822 298338 117854 298894
rect 117234 262894 117854 298338
rect 117234 262338 117266 262894
rect 117822 262338 117854 262894
rect 113514 258618 113546 259174
rect 114102 258618 114134 259174
rect 113514 223174 114134 258618
rect 116048 259174 116368 259206
rect 116048 258938 116090 259174
rect 116326 258938 116368 259174
rect 116048 258854 116368 258938
rect 116048 258618 116090 258854
rect 116326 258618 116368 258854
rect 116048 258586 116368 258618
rect 117234 226894 117854 262338
rect 117234 226338 117266 226894
rect 117822 226338 117854 226894
rect 113514 222618 113546 223174
rect 114102 222618 114134 223174
rect 113514 187174 114134 222618
rect 116048 223174 116368 223206
rect 116048 222938 116090 223174
rect 116326 222938 116368 223174
rect 116048 222854 116368 222938
rect 116048 222618 116090 222854
rect 116326 222618 116368 222854
rect 116048 222586 116368 222618
rect 117234 190894 117854 226338
rect 117234 190338 117266 190894
rect 117822 190338 117854 190894
rect 113514 186618 113546 187174
rect 114102 186618 114134 187174
rect 113514 151174 114134 186618
rect 116048 187174 116368 187206
rect 116048 186938 116090 187174
rect 116326 186938 116368 187174
rect 116048 186854 116368 186938
rect 116048 186618 116090 186854
rect 116326 186618 116368 186854
rect 116048 186586 116368 186618
rect 117234 154894 117854 190338
rect 117234 154338 117266 154894
rect 117822 154338 117854 154894
rect 113514 150618 113546 151174
rect 114102 150618 114134 151174
rect 113514 146817 114134 150618
rect 116048 151174 116368 151206
rect 116048 150938 116090 151174
rect 116326 150938 116368 151174
rect 116048 150854 116368 150938
rect 116048 150618 116090 150854
rect 116326 150618 116368 150854
rect 116048 150586 116368 150618
rect 117234 118894 117854 154338
rect 117234 118338 117266 118894
rect 117822 118338 117854 118894
rect 116048 115174 116368 115206
rect 116048 114938 116090 115174
rect 116326 114938 116368 115174
rect 116048 114854 116368 114938
rect 116048 114618 116090 114854
rect 116326 114618 116368 114854
rect 116048 114586 116368 114618
rect 109794 110898 109826 111454
rect 110382 110898 110414 111454
rect 99834 100938 99866 101494
rect 100422 100938 100454 101494
rect 99834 65494 100454 100938
rect 100688 94054 101008 94086
rect 100688 93818 100730 94054
rect 100966 93818 101008 94054
rect 100688 93734 101008 93818
rect 100688 93498 100730 93734
rect 100966 93498 101008 93734
rect 100688 93466 101008 93498
rect 108368 75454 108688 75486
rect 108368 75218 108410 75454
rect 108646 75218 108688 75454
rect 108368 75134 108688 75218
rect 108368 74898 108410 75134
rect 108646 74898 108688 75134
rect 108368 74866 108688 74898
rect 109794 75454 110414 110898
rect 117234 82894 117854 118338
rect 117234 82338 117266 82894
rect 117822 82338 117854 82894
rect 116048 79174 116368 79206
rect 116048 78938 116090 79174
rect 116326 78938 116368 79174
rect 116048 78854 116368 78938
rect 116048 78618 116090 78854
rect 116326 78618 116368 78854
rect 116048 78586 116368 78618
rect 109794 74898 109826 75454
rect 110382 74898 110414 75454
rect 99834 64938 99866 65494
rect 100422 64938 100454 65494
rect 99834 29494 100454 64938
rect 100688 58054 101008 58086
rect 100688 57818 100730 58054
rect 100966 57818 101008 58054
rect 100688 57734 101008 57818
rect 100688 57498 100730 57734
rect 100966 57498 101008 57734
rect 100688 57466 101008 57498
rect 108368 39454 108688 39486
rect 108368 39218 108410 39454
rect 108646 39218 108688 39454
rect 108368 39134 108688 39218
rect 108368 38898 108410 39134
rect 108646 38898 108688 39134
rect 108368 38866 108688 38898
rect 109794 39454 110414 74898
rect 117234 46894 117854 82338
rect 117234 46338 117266 46894
rect 117822 46338 117854 46894
rect 116048 43174 116368 43206
rect 116048 42938 116090 43174
rect 116326 42938 116368 43174
rect 116048 42854 116368 42938
rect 116048 42618 116090 42854
rect 116326 42618 116368 42854
rect 116048 42586 116368 42618
rect 109794 38898 109826 39454
rect 110382 38898 110414 39454
rect 99834 28938 99866 29494
rect 100422 28938 100454 29494
rect 99834 -7066 100454 28938
rect 100688 22054 101008 22086
rect 100688 21818 100730 22054
rect 100966 21818 101008 22054
rect 100688 21734 101008 21818
rect 100688 21498 100730 21734
rect 100966 21498 101008 21734
rect 100688 21466 101008 21498
rect 99834 -7622 99866 -7066
rect 100422 -7622 100454 -7066
rect 99834 -7654 100454 -7622
rect 109794 3454 110414 38898
rect 117234 10894 117854 46338
rect 117234 10338 117266 10894
rect 117822 10338 117854 10894
rect 116048 7174 116368 7206
rect 116048 6938 116090 7174
rect 116326 6938 116368 7174
rect 116048 6854 116368 6938
rect 116048 6618 116090 6854
rect 116326 6618 116368 6854
rect 116048 6586 116368 6618
rect 109794 2898 109826 3454
rect 110382 2898 110414 3454
rect 109794 -346 110414 2898
rect 109794 -902 109826 -346
rect 110382 -902 110414 -346
rect 109794 -7654 110414 -902
rect 113514 -1306 114134 3207
rect 113514 -1862 113546 -1306
rect 114102 -1862 114134 -1306
rect 113514 -7654 114134 -1862
rect 117234 -2266 117854 10338
rect 117234 -2822 117266 -2266
rect 117822 -2822 117854 -2266
rect 117234 -7654 117854 -2822
rect 120954 707718 121574 711590
rect 120954 707162 120986 707718
rect 121542 707162 121574 707718
rect 120954 698614 121574 707162
rect 120954 698058 120986 698614
rect 121542 698058 121574 698614
rect 120954 662614 121574 698058
rect 120954 662058 120986 662614
rect 121542 662058 121574 662614
rect 120954 626614 121574 662058
rect 120954 626058 120986 626614
rect 121542 626058 121574 626614
rect 120954 590614 121574 626058
rect 120954 590058 120986 590614
rect 121542 590058 121574 590614
rect 120954 554614 121574 590058
rect 120954 554058 120986 554614
rect 121542 554058 121574 554614
rect 120954 518614 121574 554058
rect 120954 518058 120986 518614
rect 121542 518058 121574 518614
rect 120954 482614 121574 518058
rect 120954 482058 120986 482614
rect 121542 482058 121574 482614
rect 120954 446614 121574 482058
rect 120954 446058 120986 446614
rect 121542 446058 121574 446614
rect 120954 410614 121574 446058
rect 120954 410058 120986 410614
rect 121542 410058 121574 410614
rect 120954 374614 121574 410058
rect 120954 374058 120986 374614
rect 121542 374058 121574 374614
rect 120954 338614 121574 374058
rect 120954 338058 120986 338614
rect 121542 338058 121574 338614
rect 120954 302614 121574 338058
rect 120954 302058 120986 302614
rect 121542 302058 121574 302614
rect 120954 266614 121574 302058
rect 124674 708678 125294 711590
rect 124674 708122 124706 708678
rect 125262 708122 125294 708678
rect 124674 666334 125294 708122
rect 124674 665778 124706 666334
rect 125262 665778 125294 666334
rect 124674 630334 125294 665778
rect 124674 629778 124706 630334
rect 125262 629778 125294 630334
rect 124674 594334 125294 629778
rect 124674 593778 124706 594334
rect 125262 593778 125294 594334
rect 124674 558334 125294 593778
rect 124674 557778 124706 558334
rect 125262 557778 125294 558334
rect 124674 522334 125294 557778
rect 124674 521778 124706 522334
rect 125262 521778 125294 522334
rect 124674 486334 125294 521778
rect 124674 485778 124706 486334
rect 125262 485778 125294 486334
rect 124674 450334 125294 485778
rect 124674 449778 124706 450334
rect 125262 449778 125294 450334
rect 124674 414334 125294 449778
rect 124674 413778 124706 414334
rect 125262 413778 125294 414334
rect 124674 378334 125294 413778
rect 124674 377778 124706 378334
rect 125262 377778 125294 378334
rect 124674 342334 125294 377778
rect 124674 341778 124706 342334
rect 125262 341778 125294 342334
rect 124674 306334 125294 341778
rect 124674 305778 124706 306334
rect 125262 305778 125294 306334
rect 123728 270334 124048 270366
rect 123728 270098 123770 270334
rect 124006 270098 124048 270334
rect 123728 270014 124048 270098
rect 123728 269778 123770 270014
rect 124006 269778 124048 270014
rect 123728 269746 124048 269778
rect 124674 270334 125294 305778
rect 124674 269778 124706 270334
rect 125262 269778 125294 270334
rect 120954 266058 120986 266614
rect 121542 266058 121574 266614
rect 120954 230614 121574 266058
rect 123728 234334 124048 234366
rect 123728 234098 123770 234334
rect 124006 234098 124048 234334
rect 123728 234014 124048 234098
rect 123728 233778 123770 234014
rect 124006 233778 124048 234014
rect 123728 233746 124048 233778
rect 124674 234334 125294 269778
rect 124674 233778 124706 234334
rect 125262 233778 125294 234334
rect 120954 230058 120986 230614
rect 121542 230058 121574 230614
rect 120954 194614 121574 230058
rect 123728 198334 124048 198366
rect 123728 198098 123770 198334
rect 124006 198098 124048 198334
rect 123728 198014 124048 198098
rect 123728 197778 123770 198014
rect 124006 197778 124048 198014
rect 123728 197746 124048 197778
rect 124674 198334 125294 233778
rect 124674 197778 124706 198334
rect 125262 197778 125294 198334
rect 120954 194058 120986 194614
rect 121542 194058 121574 194614
rect 120954 158614 121574 194058
rect 123728 162334 124048 162366
rect 123728 162098 123770 162334
rect 124006 162098 124048 162334
rect 123728 162014 124048 162098
rect 123728 161778 123770 162014
rect 124006 161778 124048 162014
rect 123728 161746 124048 161778
rect 124674 162334 125294 197778
rect 124674 161778 124706 162334
rect 125262 161778 125294 162334
rect 120954 158058 120986 158614
rect 121542 158058 121574 158614
rect 120954 122614 121574 158058
rect 123728 126334 124048 126366
rect 123728 126098 123770 126334
rect 124006 126098 124048 126334
rect 123728 126014 124048 126098
rect 123728 125778 123770 126014
rect 124006 125778 124048 126014
rect 123728 125746 124048 125778
rect 124674 126334 125294 161778
rect 124674 125778 124706 126334
rect 125262 125778 125294 126334
rect 120954 122058 120986 122614
rect 121542 122058 121574 122614
rect 120954 86614 121574 122058
rect 123728 90334 124048 90366
rect 123728 90098 123770 90334
rect 124006 90098 124048 90334
rect 123728 90014 124048 90098
rect 123728 89778 123770 90014
rect 124006 89778 124048 90014
rect 123728 89746 124048 89778
rect 124674 90334 125294 125778
rect 124674 89778 124706 90334
rect 125262 89778 125294 90334
rect 120954 86058 120986 86614
rect 121542 86058 121574 86614
rect 120954 50614 121574 86058
rect 123728 54334 124048 54366
rect 123728 54098 123770 54334
rect 124006 54098 124048 54334
rect 123728 54014 124048 54098
rect 123728 53778 123770 54014
rect 124006 53778 124048 54014
rect 123728 53746 124048 53778
rect 124674 54334 125294 89778
rect 124674 53778 124706 54334
rect 125262 53778 125294 54334
rect 120954 50058 120986 50614
rect 121542 50058 121574 50614
rect 120954 14614 121574 50058
rect 123728 18334 124048 18366
rect 123728 18098 123770 18334
rect 124006 18098 124048 18334
rect 123728 18014 124048 18098
rect 123728 17778 123770 18014
rect 124006 17778 124048 18014
rect 123728 17746 124048 17778
rect 124674 18334 125294 53778
rect 124674 17778 124706 18334
rect 125262 17778 125294 18334
rect 120954 14058 120986 14614
rect 121542 14058 121574 14614
rect 120954 -3226 121574 14058
rect 120954 -3782 120986 -3226
rect 121542 -3782 121574 -3226
rect 120954 -7654 121574 -3782
rect 124674 -4186 125294 17778
rect 124674 -4742 124706 -4186
rect 125262 -4742 125294 -4186
rect 124674 -7654 125294 -4742
rect 128394 709638 129014 711590
rect 128394 709082 128426 709638
rect 128982 709082 129014 709638
rect 128394 670054 129014 709082
rect 128394 669498 128426 670054
rect 128982 669498 129014 670054
rect 128394 634054 129014 669498
rect 128394 633498 128426 634054
rect 128982 633498 129014 634054
rect 128394 598054 129014 633498
rect 128394 597498 128426 598054
rect 128982 597498 129014 598054
rect 128394 562054 129014 597498
rect 128394 561498 128426 562054
rect 128982 561498 129014 562054
rect 128394 526054 129014 561498
rect 128394 525498 128426 526054
rect 128982 525498 129014 526054
rect 128394 490054 129014 525498
rect 128394 489498 128426 490054
rect 128982 489498 129014 490054
rect 128394 454054 129014 489498
rect 128394 453498 128426 454054
rect 128982 453498 129014 454054
rect 128394 418054 129014 453498
rect 128394 417498 128426 418054
rect 128982 417498 129014 418054
rect 128394 382054 129014 417498
rect 128394 381498 128426 382054
rect 128982 381498 129014 382054
rect 128394 346054 129014 381498
rect 128394 345498 128426 346054
rect 128982 345498 129014 346054
rect 128394 310054 129014 345498
rect 128394 309498 128426 310054
rect 128982 309498 129014 310054
rect 128394 274054 129014 309498
rect 132114 710598 132734 711590
rect 132114 710042 132146 710598
rect 132702 710042 132734 710598
rect 132114 673774 132734 710042
rect 132114 673218 132146 673774
rect 132702 673218 132734 673774
rect 132114 637774 132734 673218
rect 132114 637218 132146 637774
rect 132702 637218 132734 637774
rect 132114 601774 132734 637218
rect 132114 601218 132146 601774
rect 132702 601218 132734 601774
rect 132114 565774 132734 601218
rect 132114 565218 132146 565774
rect 132702 565218 132734 565774
rect 132114 529774 132734 565218
rect 132114 529218 132146 529774
rect 132702 529218 132734 529774
rect 132114 493774 132734 529218
rect 132114 493218 132146 493774
rect 132702 493218 132734 493774
rect 132114 457774 132734 493218
rect 132114 457218 132146 457774
rect 132702 457218 132734 457774
rect 132114 421774 132734 457218
rect 132114 421218 132146 421774
rect 132702 421218 132734 421774
rect 132114 385774 132734 421218
rect 132114 385218 132146 385774
rect 132702 385218 132734 385774
rect 132114 349774 132734 385218
rect 132114 349218 132146 349774
rect 132702 349218 132734 349774
rect 132114 313774 132734 349218
rect 132114 313218 132146 313774
rect 132702 313218 132734 313774
rect 132114 277774 132734 313218
rect 132114 277218 132146 277774
rect 132702 277218 132734 277774
rect 128394 273498 128426 274054
rect 128982 273498 129014 274054
rect 128394 238054 129014 273498
rect 131408 274054 131728 274086
rect 131408 273818 131450 274054
rect 131686 273818 131728 274054
rect 131408 273734 131728 273818
rect 131408 273498 131450 273734
rect 131686 273498 131728 273734
rect 131408 273466 131728 273498
rect 132114 241774 132734 277218
rect 132114 241218 132146 241774
rect 132702 241218 132734 241774
rect 128394 237498 128426 238054
rect 128982 237498 129014 238054
rect 128394 202054 129014 237498
rect 131408 238054 131728 238086
rect 131408 237818 131450 238054
rect 131686 237818 131728 238054
rect 131408 237734 131728 237818
rect 131408 237498 131450 237734
rect 131686 237498 131728 237734
rect 131408 237466 131728 237498
rect 132114 205774 132734 241218
rect 132114 205218 132146 205774
rect 132702 205218 132734 205774
rect 128394 201498 128426 202054
rect 128982 201498 129014 202054
rect 128394 166054 129014 201498
rect 131408 202054 131728 202086
rect 131408 201818 131450 202054
rect 131686 201818 131728 202054
rect 131408 201734 131728 201818
rect 131408 201498 131450 201734
rect 131686 201498 131728 201734
rect 131408 201466 131728 201498
rect 132114 169774 132734 205218
rect 132114 169218 132146 169774
rect 132702 169218 132734 169774
rect 128394 165498 128426 166054
rect 128982 165498 129014 166054
rect 128394 130054 129014 165498
rect 131408 166054 131728 166086
rect 131408 165818 131450 166054
rect 131686 165818 131728 166054
rect 131408 165734 131728 165818
rect 131408 165498 131450 165734
rect 131686 165498 131728 165734
rect 131408 165466 131728 165498
rect 132114 133774 132734 169218
rect 132114 133218 132146 133774
rect 132702 133218 132734 133774
rect 128394 129498 128426 130054
rect 128982 129498 129014 130054
rect 128394 94054 129014 129498
rect 131408 130054 131728 130086
rect 131408 129818 131450 130054
rect 131686 129818 131728 130054
rect 131408 129734 131728 129818
rect 131408 129498 131450 129734
rect 131686 129498 131728 129734
rect 131408 129466 131728 129498
rect 132114 97774 132734 133218
rect 132114 97218 132146 97774
rect 132702 97218 132734 97774
rect 128394 93498 128426 94054
rect 128982 93498 129014 94054
rect 128394 58054 129014 93498
rect 131408 94054 131728 94086
rect 131408 93818 131450 94054
rect 131686 93818 131728 94054
rect 131408 93734 131728 93818
rect 131408 93498 131450 93734
rect 131686 93498 131728 93734
rect 131408 93466 131728 93498
rect 132114 61774 132734 97218
rect 132114 61218 132146 61774
rect 132702 61218 132734 61774
rect 128394 57498 128426 58054
rect 128982 57498 129014 58054
rect 128394 22054 129014 57498
rect 131408 58054 131728 58086
rect 131408 57818 131450 58054
rect 131686 57818 131728 58054
rect 131408 57734 131728 57818
rect 131408 57498 131450 57734
rect 131686 57498 131728 57734
rect 131408 57466 131728 57498
rect 132114 25774 132734 61218
rect 132114 25218 132146 25774
rect 132702 25218 132734 25774
rect 128394 21498 128426 22054
rect 128982 21498 129014 22054
rect 128394 -5146 129014 21498
rect 131408 22054 131728 22086
rect 131408 21818 131450 22054
rect 131686 21818 131728 22054
rect 131408 21734 131728 21818
rect 131408 21498 131450 21734
rect 131686 21498 131728 21734
rect 131408 21466 131728 21498
rect 128394 -5702 128426 -5146
rect 128982 -5702 129014 -5146
rect 128394 -7654 129014 -5702
rect 132114 -6106 132734 25218
rect 132114 -6662 132146 -6106
rect 132702 -6662 132734 -6106
rect 132114 -7654 132734 -6662
rect 135834 711558 136454 711590
rect 135834 711002 135866 711558
rect 136422 711002 136454 711558
rect 135834 677494 136454 711002
rect 135834 676938 135866 677494
rect 136422 676938 136454 677494
rect 135834 641494 136454 676938
rect 135834 640938 135866 641494
rect 136422 640938 136454 641494
rect 135834 605494 136454 640938
rect 135834 604938 135866 605494
rect 136422 604938 136454 605494
rect 135834 569494 136454 604938
rect 135834 568938 135866 569494
rect 136422 568938 136454 569494
rect 135834 533494 136454 568938
rect 135834 532938 135866 533494
rect 136422 532938 136454 533494
rect 135834 497494 136454 532938
rect 135834 496938 135866 497494
rect 136422 496938 136454 497494
rect 135834 461494 136454 496938
rect 135834 460938 135866 461494
rect 136422 460938 136454 461494
rect 135834 425494 136454 460938
rect 135834 424938 135866 425494
rect 136422 424938 136454 425494
rect 135834 389494 136454 424938
rect 135834 388938 135866 389494
rect 136422 388938 136454 389494
rect 135834 353494 136454 388938
rect 135834 352938 135866 353494
rect 136422 352938 136454 353494
rect 135834 317494 136454 352938
rect 135834 316938 135866 317494
rect 136422 316938 136454 317494
rect 135834 281494 136454 316938
rect 135834 280938 135866 281494
rect 136422 280938 136454 281494
rect 135834 245494 136454 280938
rect 145794 704838 146414 711590
rect 145794 704282 145826 704838
rect 146382 704282 146414 704838
rect 145794 687454 146414 704282
rect 145794 686898 145826 687454
rect 146382 686898 146414 687454
rect 145794 651454 146414 686898
rect 145794 650898 145826 651454
rect 146382 650898 146414 651454
rect 145794 615454 146414 650898
rect 145794 614898 145826 615454
rect 146382 614898 146414 615454
rect 145794 579454 146414 614898
rect 145794 578898 145826 579454
rect 146382 578898 146414 579454
rect 145794 543454 146414 578898
rect 145794 542898 145826 543454
rect 146382 542898 146414 543454
rect 145794 507454 146414 542898
rect 145794 506898 145826 507454
rect 146382 506898 146414 507454
rect 145794 471454 146414 506898
rect 145794 470898 145826 471454
rect 146382 470898 146414 471454
rect 145794 435454 146414 470898
rect 145794 434898 145826 435454
rect 146382 434898 146414 435454
rect 145794 399454 146414 434898
rect 145794 398898 145826 399454
rect 146382 398898 146414 399454
rect 145794 363454 146414 398898
rect 145794 362898 145826 363454
rect 146382 362898 146414 363454
rect 145794 327454 146414 362898
rect 145794 326898 145826 327454
rect 146382 326898 146414 327454
rect 145794 291454 146414 326898
rect 145794 290898 145826 291454
rect 146382 290898 146414 291454
rect 139088 255454 139408 255486
rect 139088 255218 139130 255454
rect 139366 255218 139408 255454
rect 139088 255134 139408 255218
rect 139088 254898 139130 255134
rect 139366 254898 139408 255134
rect 139088 254866 139408 254898
rect 145794 255454 146414 290898
rect 149514 705798 150134 711590
rect 149514 705242 149546 705798
rect 150102 705242 150134 705798
rect 149514 691174 150134 705242
rect 149514 690618 149546 691174
rect 150102 690618 150134 691174
rect 149514 655174 150134 690618
rect 149514 654618 149546 655174
rect 150102 654618 150134 655174
rect 149514 619174 150134 654618
rect 149514 618618 149546 619174
rect 150102 618618 150134 619174
rect 149514 583174 150134 618618
rect 149514 582618 149546 583174
rect 150102 582618 150134 583174
rect 149514 547174 150134 582618
rect 149514 546618 149546 547174
rect 150102 546618 150134 547174
rect 149514 511174 150134 546618
rect 149514 510618 149546 511174
rect 150102 510618 150134 511174
rect 149514 475174 150134 510618
rect 149514 474618 149546 475174
rect 150102 474618 150134 475174
rect 149514 439174 150134 474618
rect 149514 438618 149546 439174
rect 150102 438618 150134 439174
rect 149514 403174 150134 438618
rect 149514 402618 149546 403174
rect 150102 402618 150134 403174
rect 149514 367174 150134 402618
rect 149514 366618 149546 367174
rect 150102 366618 150134 367174
rect 149514 331174 150134 366618
rect 149514 330618 149546 331174
rect 150102 330618 150134 331174
rect 149514 295174 150134 330618
rect 149514 294618 149546 295174
rect 150102 294618 150134 295174
rect 146768 259174 147088 259206
rect 146768 258938 146810 259174
rect 147046 258938 147088 259174
rect 146768 258854 147088 258938
rect 146768 258618 146810 258854
rect 147046 258618 147088 258854
rect 146768 258586 147088 258618
rect 149514 259174 150134 294618
rect 149514 258618 149546 259174
rect 150102 258618 150134 259174
rect 145794 254898 145826 255454
rect 146382 254898 146414 255454
rect 135834 244938 135866 245494
rect 136422 244938 136454 245494
rect 135834 209494 136454 244938
rect 139088 219454 139408 219486
rect 139088 219218 139130 219454
rect 139366 219218 139408 219454
rect 139088 219134 139408 219218
rect 139088 218898 139130 219134
rect 139366 218898 139408 219134
rect 139088 218866 139408 218898
rect 145794 219454 146414 254898
rect 146768 223174 147088 223206
rect 146768 222938 146810 223174
rect 147046 222938 147088 223174
rect 146768 222854 147088 222938
rect 146768 222618 146810 222854
rect 147046 222618 147088 222854
rect 146768 222586 147088 222618
rect 149514 223174 150134 258618
rect 149514 222618 149546 223174
rect 150102 222618 150134 223174
rect 145794 218898 145826 219454
rect 146382 218898 146414 219454
rect 135834 208938 135866 209494
rect 136422 208938 136454 209494
rect 135834 173494 136454 208938
rect 139088 183454 139408 183486
rect 139088 183218 139130 183454
rect 139366 183218 139408 183454
rect 139088 183134 139408 183218
rect 139088 182898 139130 183134
rect 139366 182898 139408 183134
rect 139088 182866 139408 182898
rect 145794 183454 146414 218898
rect 146768 187174 147088 187206
rect 146768 186938 146810 187174
rect 147046 186938 147088 187174
rect 146768 186854 147088 186938
rect 146768 186618 146810 186854
rect 147046 186618 147088 186854
rect 146768 186586 147088 186618
rect 149514 187174 150134 222618
rect 149514 186618 149546 187174
rect 150102 186618 150134 187174
rect 145794 182898 145826 183454
rect 146382 182898 146414 183454
rect 135834 172938 135866 173494
rect 136422 172938 136454 173494
rect 135834 137494 136454 172938
rect 139088 147454 139408 147486
rect 139088 147218 139130 147454
rect 139366 147218 139408 147454
rect 139088 147134 139408 147218
rect 139088 146898 139130 147134
rect 139366 146898 139408 147134
rect 139088 146866 139408 146898
rect 145794 147454 146414 182898
rect 146768 151174 147088 151206
rect 146768 150938 146810 151174
rect 147046 150938 147088 151174
rect 146768 150854 147088 150938
rect 146768 150618 146810 150854
rect 147046 150618 147088 150854
rect 146768 150586 147088 150618
rect 149514 151174 150134 186618
rect 149514 150618 149546 151174
rect 150102 150618 150134 151174
rect 145794 146898 145826 147454
rect 146382 146898 146414 147454
rect 135834 136938 135866 137494
rect 136422 136938 136454 137494
rect 135834 101494 136454 136938
rect 139088 111454 139408 111486
rect 139088 111218 139130 111454
rect 139366 111218 139408 111454
rect 139088 111134 139408 111218
rect 139088 110898 139130 111134
rect 139366 110898 139408 111134
rect 139088 110866 139408 110898
rect 145794 111454 146414 146898
rect 146768 115174 147088 115206
rect 146768 114938 146810 115174
rect 147046 114938 147088 115174
rect 146768 114854 147088 114938
rect 146768 114618 146810 114854
rect 147046 114618 147088 114854
rect 146768 114586 147088 114618
rect 149514 115174 150134 150618
rect 149514 114618 149546 115174
rect 150102 114618 150134 115174
rect 145794 110898 145826 111454
rect 146382 110898 146414 111454
rect 135834 100938 135866 101494
rect 136422 100938 136454 101494
rect 135834 65494 136454 100938
rect 139088 75454 139408 75486
rect 139088 75218 139130 75454
rect 139366 75218 139408 75454
rect 139088 75134 139408 75218
rect 139088 74898 139130 75134
rect 139366 74898 139408 75134
rect 139088 74866 139408 74898
rect 145794 75454 146414 110898
rect 146768 79174 147088 79206
rect 146768 78938 146810 79174
rect 147046 78938 147088 79174
rect 146768 78854 147088 78938
rect 146768 78618 146810 78854
rect 147046 78618 147088 78854
rect 146768 78586 147088 78618
rect 149514 79174 150134 114618
rect 149514 78618 149546 79174
rect 150102 78618 150134 79174
rect 145794 74898 145826 75454
rect 146382 74898 146414 75454
rect 135834 64938 135866 65494
rect 136422 64938 136454 65494
rect 135834 29494 136454 64938
rect 139088 39454 139408 39486
rect 139088 39218 139130 39454
rect 139366 39218 139408 39454
rect 139088 39134 139408 39218
rect 139088 38898 139130 39134
rect 139366 38898 139408 39134
rect 139088 38866 139408 38898
rect 145794 39454 146414 74898
rect 146768 43174 147088 43206
rect 146768 42938 146810 43174
rect 147046 42938 147088 43174
rect 146768 42854 147088 42938
rect 146768 42618 146810 42854
rect 147046 42618 147088 42854
rect 146768 42586 147088 42618
rect 149514 43174 150134 78618
rect 149514 42618 149546 43174
rect 150102 42618 150134 43174
rect 145794 38898 145826 39454
rect 146382 38898 146414 39454
rect 135834 28938 135866 29494
rect 136422 28938 136454 29494
rect 135834 -7066 136454 28938
rect 135834 -7622 135866 -7066
rect 136422 -7622 136454 -7066
rect 135834 -7654 136454 -7622
rect 145794 3454 146414 38898
rect 146768 7174 147088 7206
rect 146768 6938 146810 7174
rect 147046 6938 147088 7174
rect 146768 6854 147088 6938
rect 146768 6618 146810 6854
rect 147046 6618 147088 6854
rect 146768 6586 147088 6618
rect 149514 7174 150134 42618
rect 149514 6618 149546 7174
rect 150102 6618 150134 7174
rect 145794 2898 145826 3454
rect 146382 2898 146414 3454
rect 145794 -346 146414 2898
rect 145794 -902 145826 -346
rect 146382 -902 146414 -346
rect 145794 -7654 146414 -902
rect 149514 -1306 150134 6618
rect 149514 -1862 149546 -1306
rect 150102 -1862 150134 -1306
rect 149514 -7654 150134 -1862
rect 153234 706758 153854 711590
rect 153234 706202 153266 706758
rect 153822 706202 153854 706758
rect 153234 694894 153854 706202
rect 153234 694338 153266 694894
rect 153822 694338 153854 694894
rect 153234 658894 153854 694338
rect 153234 658338 153266 658894
rect 153822 658338 153854 658894
rect 153234 622894 153854 658338
rect 153234 622338 153266 622894
rect 153822 622338 153854 622894
rect 153234 586894 153854 622338
rect 153234 586338 153266 586894
rect 153822 586338 153854 586894
rect 153234 550894 153854 586338
rect 153234 550338 153266 550894
rect 153822 550338 153854 550894
rect 153234 514894 153854 550338
rect 153234 514338 153266 514894
rect 153822 514338 153854 514894
rect 153234 478894 153854 514338
rect 153234 478338 153266 478894
rect 153822 478338 153854 478894
rect 153234 442894 153854 478338
rect 153234 442338 153266 442894
rect 153822 442338 153854 442894
rect 153234 406894 153854 442338
rect 153234 406338 153266 406894
rect 153822 406338 153854 406894
rect 153234 370894 153854 406338
rect 153234 370338 153266 370894
rect 153822 370338 153854 370894
rect 153234 334894 153854 370338
rect 153234 334338 153266 334894
rect 153822 334338 153854 334894
rect 153234 298894 153854 334338
rect 153234 298338 153266 298894
rect 153822 298338 153854 298894
rect 153234 262894 153854 298338
rect 156954 707718 157574 711590
rect 156954 707162 156986 707718
rect 157542 707162 157574 707718
rect 156954 698614 157574 707162
rect 156954 698058 156986 698614
rect 157542 698058 157574 698614
rect 156954 662614 157574 698058
rect 156954 662058 156986 662614
rect 157542 662058 157574 662614
rect 156954 626614 157574 662058
rect 156954 626058 156986 626614
rect 157542 626058 157574 626614
rect 156954 590614 157574 626058
rect 156954 590058 156986 590614
rect 157542 590058 157574 590614
rect 156954 554614 157574 590058
rect 156954 554058 156986 554614
rect 157542 554058 157574 554614
rect 156954 518614 157574 554058
rect 156954 518058 156986 518614
rect 157542 518058 157574 518614
rect 156954 482614 157574 518058
rect 156954 482058 156986 482614
rect 157542 482058 157574 482614
rect 156954 446614 157574 482058
rect 156954 446058 156986 446614
rect 157542 446058 157574 446614
rect 156954 410614 157574 446058
rect 156954 410058 156986 410614
rect 157542 410058 157574 410614
rect 156954 374614 157574 410058
rect 156954 374058 156986 374614
rect 157542 374058 157574 374614
rect 156954 338614 157574 374058
rect 156954 338058 156986 338614
rect 157542 338058 157574 338614
rect 156954 302614 157574 338058
rect 156954 302058 156986 302614
rect 157542 302058 157574 302614
rect 154448 270334 154768 270366
rect 154448 270098 154490 270334
rect 154726 270098 154768 270334
rect 154448 270014 154768 270098
rect 154448 269778 154490 270014
rect 154726 269778 154768 270014
rect 154448 269746 154768 269778
rect 153234 262338 153266 262894
rect 153822 262338 153854 262894
rect 153234 226894 153854 262338
rect 156954 266614 157574 302058
rect 156954 266058 156986 266614
rect 157542 266058 157574 266614
rect 154448 234334 154768 234366
rect 154448 234098 154490 234334
rect 154726 234098 154768 234334
rect 154448 234014 154768 234098
rect 154448 233778 154490 234014
rect 154726 233778 154768 234014
rect 154448 233746 154768 233778
rect 153234 226338 153266 226894
rect 153822 226338 153854 226894
rect 153234 190894 153854 226338
rect 156954 230614 157574 266058
rect 156954 230058 156986 230614
rect 157542 230058 157574 230614
rect 154448 198334 154768 198366
rect 154448 198098 154490 198334
rect 154726 198098 154768 198334
rect 154448 198014 154768 198098
rect 154448 197778 154490 198014
rect 154726 197778 154768 198014
rect 154448 197746 154768 197778
rect 153234 190338 153266 190894
rect 153822 190338 153854 190894
rect 153234 154894 153854 190338
rect 156954 194614 157574 230058
rect 156954 194058 156986 194614
rect 157542 194058 157574 194614
rect 154448 162334 154768 162366
rect 154448 162098 154490 162334
rect 154726 162098 154768 162334
rect 154448 162014 154768 162098
rect 154448 161778 154490 162014
rect 154726 161778 154768 162014
rect 154448 161746 154768 161778
rect 153234 154338 153266 154894
rect 153822 154338 153854 154894
rect 153234 118894 153854 154338
rect 156954 158614 157574 194058
rect 156954 158058 156986 158614
rect 157542 158058 157574 158614
rect 154448 126334 154768 126366
rect 154448 126098 154490 126334
rect 154726 126098 154768 126334
rect 154448 126014 154768 126098
rect 154448 125778 154490 126014
rect 154726 125778 154768 126014
rect 154448 125746 154768 125778
rect 153234 118338 153266 118894
rect 153822 118338 153854 118894
rect 153234 82894 153854 118338
rect 156954 122614 157574 158058
rect 156954 122058 156986 122614
rect 157542 122058 157574 122614
rect 154448 90334 154768 90366
rect 154448 90098 154490 90334
rect 154726 90098 154768 90334
rect 154448 90014 154768 90098
rect 154448 89778 154490 90014
rect 154726 89778 154768 90014
rect 154448 89746 154768 89778
rect 153234 82338 153266 82894
rect 153822 82338 153854 82894
rect 153234 46894 153854 82338
rect 156954 86614 157574 122058
rect 156954 86058 156986 86614
rect 157542 86058 157574 86614
rect 154448 54334 154768 54366
rect 154448 54098 154490 54334
rect 154726 54098 154768 54334
rect 154448 54014 154768 54098
rect 154448 53778 154490 54014
rect 154726 53778 154768 54014
rect 154448 53746 154768 53778
rect 153234 46338 153266 46894
rect 153822 46338 153854 46894
rect 153234 10894 153854 46338
rect 156954 50614 157574 86058
rect 156954 50058 156986 50614
rect 157542 50058 157574 50614
rect 154448 18334 154768 18366
rect 154448 18098 154490 18334
rect 154726 18098 154768 18334
rect 154448 18014 154768 18098
rect 154448 17778 154490 18014
rect 154726 17778 154768 18014
rect 154448 17746 154768 17778
rect 153234 10338 153266 10894
rect 153822 10338 153854 10894
rect 153234 -2266 153854 10338
rect 153234 -2822 153266 -2266
rect 153822 -2822 153854 -2266
rect 153234 -7654 153854 -2822
rect 156954 14614 157574 50058
rect 156954 14058 156986 14614
rect 157542 14058 157574 14614
rect 156954 -3226 157574 14058
rect 156954 -3782 156986 -3226
rect 157542 -3782 157574 -3226
rect 156954 -7654 157574 -3782
rect 160674 708678 161294 711590
rect 160674 708122 160706 708678
rect 161262 708122 161294 708678
rect 160674 666334 161294 708122
rect 160674 665778 160706 666334
rect 161262 665778 161294 666334
rect 160674 630334 161294 665778
rect 160674 629778 160706 630334
rect 161262 629778 161294 630334
rect 160674 594334 161294 629778
rect 160674 593778 160706 594334
rect 161262 593778 161294 594334
rect 160674 558334 161294 593778
rect 160674 557778 160706 558334
rect 161262 557778 161294 558334
rect 160674 522334 161294 557778
rect 160674 521778 160706 522334
rect 161262 521778 161294 522334
rect 160674 486334 161294 521778
rect 160674 485778 160706 486334
rect 161262 485778 161294 486334
rect 160674 450334 161294 485778
rect 160674 449778 160706 450334
rect 161262 449778 161294 450334
rect 160674 414334 161294 449778
rect 160674 413778 160706 414334
rect 161262 413778 161294 414334
rect 160674 378334 161294 413778
rect 160674 377778 160706 378334
rect 161262 377778 161294 378334
rect 160674 342334 161294 377778
rect 160674 341778 160706 342334
rect 161262 341778 161294 342334
rect 160674 306334 161294 341778
rect 160674 305778 160706 306334
rect 161262 305778 161294 306334
rect 160674 270334 161294 305778
rect 164394 709638 165014 711590
rect 164394 709082 164426 709638
rect 164982 709082 165014 709638
rect 164394 670054 165014 709082
rect 164394 669498 164426 670054
rect 164982 669498 165014 670054
rect 164394 634054 165014 669498
rect 164394 633498 164426 634054
rect 164982 633498 165014 634054
rect 164394 598054 165014 633498
rect 164394 597498 164426 598054
rect 164982 597498 165014 598054
rect 164394 562054 165014 597498
rect 164394 561498 164426 562054
rect 164982 561498 165014 562054
rect 164394 526054 165014 561498
rect 164394 525498 164426 526054
rect 164982 525498 165014 526054
rect 164394 490054 165014 525498
rect 164394 489498 164426 490054
rect 164982 489498 165014 490054
rect 164394 454054 165014 489498
rect 164394 453498 164426 454054
rect 164982 453498 165014 454054
rect 164394 418054 165014 453498
rect 164394 417498 164426 418054
rect 164982 417498 165014 418054
rect 164394 382054 165014 417498
rect 164394 381498 164426 382054
rect 164982 381498 165014 382054
rect 164394 346054 165014 381498
rect 164394 345498 164426 346054
rect 164982 345498 165014 346054
rect 164394 310054 165014 345498
rect 164394 309498 164426 310054
rect 164982 309498 165014 310054
rect 162128 274054 162448 274086
rect 162128 273818 162170 274054
rect 162406 273818 162448 274054
rect 162128 273734 162448 273818
rect 162128 273498 162170 273734
rect 162406 273498 162448 273734
rect 162128 273466 162448 273498
rect 164394 274054 165014 309498
rect 164394 273498 164426 274054
rect 164982 273498 165014 274054
rect 160674 269778 160706 270334
rect 161262 269778 161294 270334
rect 160674 234334 161294 269778
rect 162128 238054 162448 238086
rect 162128 237818 162170 238054
rect 162406 237818 162448 238054
rect 162128 237734 162448 237818
rect 162128 237498 162170 237734
rect 162406 237498 162448 237734
rect 162128 237466 162448 237498
rect 164394 238054 165014 273498
rect 164394 237498 164426 238054
rect 164982 237498 165014 238054
rect 160674 233778 160706 234334
rect 161262 233778 161294 234334
rect 160674 198334 161294 233778
rect 162128 202054 162448 202086
rect 162128 201818 162170 202054
rect 162406 201818 162448 202054
rect 162128 201734 162448 201818
rect 162128 201498 162170 201734
rect 162406 201498 162448 201734
rect 162128 201466 162448 201498
rect 164394 202054 165014 237498
rect 164394 201498 164426 202054
rect 164982 201498 165014 202054
rect 160674 197778 160706 198334
rect 161262 197778 161294 198334
rect 160674 162334 161294 197778
rect 162128 166054 162448 166086
rect 162128 165818 162170 166054
rect 162406 165818 162448 166054
rect 162128 165734 162448 165818
rect 162128 165498 162170 165734
rect 162406 165498 162448 165734
rect 162128 165466 162448 165498
rect 164394 166054 165014 201498
rect 164394 165498 164426 166054
rect 164982 165498 165014 166054
rect 160674 161778 160706 162334
rect 161262 161778 161294 162334
rect 160674 126334 161294 161778
rect 162128 130054 162448 130086
rect 162128 129818 162170 130054
rect 162406 129818 162448 130054
rect 162128 129734 162448 129818
rect 162128 129498 162170 129734
rect 162406 129498 162448 129734
rect 162128 129466 162448 129498
rect 164394 130054 165014 165498
rect 164394 129498 164426 130054
rect 164982 129498 165014 130054
rect 160674 125778 160706 126334
rect 161262 125778 161294 126334
rect 160674 90334 161294 125778
rect 162128 94054 162448 94086
rect 162128 93818 162170 94054
rect 162406 93818 162448 94054
rect 162128 93734 162448 93818
rect 162128 93498 162170 93734
rect 162406 93498 162448 93734
rect 162128 93466 162448 93498
rect 164394 94054 165014 129498
rect 164394 93498 164426 94054
rect 164982 93498 165014 94054
rect 160674 89778 160706 90334
rect 161262 89778 161294 90334
rect 160674 54334 161294 89778
rect 162128 58054 162448 58086
rect 162128 57818 162170 58054
rect 162406 57818 162448 58054
rect 162128 57734 162448 57818
rect 162128 57498 162170 57734
rect 162406 57498 162448 57734
rect 162128 57466 162448 57498
rect 164394 58054 165014 93498
rect 164394 57498 164426 58054
rect 164982 57498 165014 58054
rect 160674 53778 160706 54334
rect 161262 53778 161294 54334
rect 160674 18334 161294 53778
rect 162128 22054 162448 22086
rect 162128 21818 162170 22054
rect 162406 21818 162448 22054
rect 162128 21734 162448 21818
rect 162128 21498 162170 21734
rect 162406 21498 162448 21734
rect 162128 21466 162448 21498
rect 164394 22054 165014 57498
rect 164394 21498 164426 22054
rect 164982 21498 165014 22054
rect 160674 17778 160706 18334
rect 161262 17778 161294 18334
rect 160674 -4186 161294 17778
rect 160674 -4742 160706 -4186
rect 161262 -4742 161294 -4186
rect 160674 -7654 161294 -4742
rect 164394 -5146 165014 21498
rect 164394 -5702 164426 -5146
rect 164982 -5702 165014 -5146
rect 164394 -7654 165014 -5702
rect 168114 710598 168734 711590
rect 168114 710042 168146 710598
rect 168702 710042 168734 710598
rect 168114 673774 168734 710042
rect 168114 673218 168146 673774
rect 168702 673218 168734 673774
rect 168114 637774 168734 673218
rect 168114 637218 168146 637774
rect 168702 637218 168734 637774
rect 168114 601774 168734 637218
rect 168114 601218 168146 601774
rect 168702 601218 168734 601774
rect 168114 565774 168734 601218
rect 168114 565218 168146 565774
rect 168702 565218 168734 565774
rect 168114 529774 168734 565218
rect 168114 529218 168146 529774
rect 168702 529218 168734 529774
rect 168114 493774 168734 529218
rect 168114 493218 168146 493774
rect 168702 493218 168734 493774
rect 168114 457774 168734 493218
rect 168114 457218 168146 457774
rect 168702 457218 168734 457774
rect 168114 421774 168734 457218
rect 168114 421218 168146 421774
rect 168702 421218 168734 421774
rect 168114 385774 168734 421218
rect 168114 385218 168146 385774
rect 168702 385218 168734 385774
rect 168114 349774 168734 385218
rect 168114 349218 168146 349774
rect 168702 349218 168734 349774
rect 168114 313774 168734 349218
rect 168114 313218 168146 313774
rect 168702 313218 168734 313774
rect 168114 277774 168734 313218
rect 168114 277218 168146 277774
rect 168702 277218 168734 277774
rect 168114 241774 168734 277218
rect 171834 711558 172454 711590
rect 171834 711002 171866 711558
rect 172422 711002 172454 711558
rect 171834 677494 172454 711002
rect 171834 676938 171866 677494
rect 172422 676938 172454 677494
rect 171834 641494 172454 676938
rect 171834 640938 171866 641494
rect 172422 640938 172454 641494
rect 171834 605494 172454 640938
rect 171834 604938 171866 605494
rect 172422 604938 172454 605494
rect 171834 569494 172454 604938
rect 171834 568938 171866 569494
rect 172422 568938 172454 569494
rect 171834 533494 172454 568938
rect 171834 532938 171866 533494
rect 172422 532938 172454 533494
rect 171834 497494 172454 532938
rect 171834 496938 171866 497494
rect 172422 496938 172454 497494
rect 171834 461494 172454 496938
rect 171834 460938 171866 461494
rect 172422 460938 172454 461494
rect 171834 425494 172454 460938
rect 171834 424938 171866 425494
rect 172422 424938 172454 425494
rect 171834 389494 172454 424938
rect 171834 388938 171866 389494
rect 172422 388938 172454 389494
rect 171834 353494 172454 388938
rect 171834 352938 171866 353494
rect 172422 352938 172454 353494
rect 171834 317494 172454 352938
rect 171834 316938 171866 317494
rect 172422 316938 172454 317494
rect 171834 281494 172454 316938
rect 171834 280938 171866 281494
rect 172422 280938 172454 281494
rect 169808 255454 170128 255486
rect 169808 255218 169850 255454
rect 170086 255218 170128 255454
rect 169808 255134 170128 255218
rect 169808 254898 169850 255134
rect 170086 254898 170128 255134
rect 169808 254866 170128 254898
rect 168114 241218 168146 241774
rect 168702 241218 168734 241774
rect 168114 205774 168734 241218
rect 171834 245494 172454 280938
rect 181794 704838 182414 711590
rect 181794 704282 181826 704838
rect 182382 704282 182414 704838
rect 181794 687454 182414 704282
rect 181794 686898 181826 687454
rect 182382 686898 182414 687454
rect 181794 651454 182414 686898
rect 181794 650898 181826 651454
rect 182382 650898 182414 651454
rect 181794 615454 182414 650898
rect 181794 614898 181826 615454
rect 182382 614898 182414 615454
rect 181794 579454 182414 614898
rect 181794 578898 181826 579454
rect 182382 578898 182414 579454
rect 181794 543454 182414 578898
rect 181794 542898 181826 543454
rect 182382 542898 182414 543454
rect 181794 507454 182414 542898
rect 181794 506898 181826 507454
rect 182382 506898 182414 507454
rect 181794 471454 182414 506898
rect 181794 470898 181826 471454
rect 182382 470898 182414 471454
rect 181794 435454 182414 470898
rect 181794 434898 181826 435454
rect 182382 434898 182414 435454
rect 181794 399454 182414 434898
rect 181794 398898 181826 399454
rect 182382 398898 182414 399454
rect 181794 363454 182414 398898
rect 181794 362898 181826 363454
rect 182382 362898 182414 363454
rect 181794 327454 182414 362898
rect 181794 326898 181826 327454
rect 182382 326898 182414 327454
rect 181794 291454 182414 326898
rect 181794 290898 181826 291454
rect 182382 290898 182414 291454
rect 177488 259174 177808 259206
rect 177488 258938 177530 259174
rect 177766 258938 177808 259174
rect 177488 258854 177808 258938
rect 177488 258618 177530 258854
rect 177766 258618 177808 258854
rect 177488 258586 177808 258618
rect 171834 244938 171866 245494
rect 172422 244938 172454 245494
rect 169808 219454 170128 219486
rect 169808 219218 169850 219454
rect 170086 219218 170128 219454
rect 169808 219134 170128 219218
rect 169808 218898 169850 219134
rect 170086 218898 170128 219134
rect 169808 218866 170128 218898
rect 168114 205218 168146 205774
rect 168702 205218 168734 205774
rect 168114 169774 168734 205218
rect 171834 209494 172454 244938
rect 181794 255454 182414 290898
rect 185514 705798 186134 711590
rect 185514 705242 185546 705798
rect 186102 705242 186134 705798
rect 185514 691174 186134 705242
rect 185514 690618 185546 691174
rect 186102 690618 186134 691174
rect 185514 655174 186134 690618
rect 185514 654618 185546 655174
rect 186102 654618 186134 655174
rect 185514 619174 186134 654618
rect 185514 618618 185546 619174
rect 186102 618618 186134 619174
rect 185514 583174 186134 618618
rect 185514 582618 185546 583174
rect 186102 582618 186134 583174
rect 185514 547174 186134 582618
rect 185514 546618 185546 547174
rect 186102 546618 186134 547174
rect 185514 511174 186134 546618
rect 185514 510618 185546 511174
rect 186102 510618 186134 511174
rect 185514 475174 186134 510618
rect 185514 474618 185546 475174
rect 186102 474618 186134 475174
rect 185514 439174 186134 474618
rect 185514 438618 185546 439174
rect 186102 438618 186134 439174
rect 185514 403174 186134 438618
rect 185514 402618 185546 403174
rect 186102 402618 186134 403174
rect 185514 367174 186134 402618
rect 185514 366618 185546 367174
rect 186102 366618 186134 367174
rect 185514 331174 186134 366618
rect 185514 330618 185546 331174
rect 186102 330618 186134 331174
rect 185514 295174 186134 330618
rect 185514 294618 185546 295174
rect 186102 294618 186134 295174
rect 185514 282628 186134 294618
rect 189234 706758 189854 711590
rect 189234 706202 189266 706758
rect 189822 706202 189854 706758
rect 189234 694894 189854 706202
rect 189234 694338 189266 694894
rect 189822 694338 189854 694894
rect 189234 658894 189854 694338
rect 189234 658338 189266 658894
rect 189822 658338 189854 658894
rect 189234 622894 189854 658338
rect 189234 622338 189266 622894
rect 189822 622338 189854 622894
rect 189234 586894 189854 622338
rect 189234 586338 189266 586894
rect 189822 586338 189854 586894
rect 189234 550894 189854 586338
rect 189234 550338 189266 550894
rect 189822 550338 189854 550894
rect 189234 514894 189854 550338
rect 189234 514338 189266 514894
rect 189822 514338 189854 514894
rect 189234 478894 189854 514338
rect 189234 478338 189266 478894
rect 189822 478338 189854 478894
rect 189234 442894 189854 478338
rect 189234 442338 189266 442894
rect 189822 442338 189854 442894
rect 189234 406894 189854 442338
rect 189234 406338 189266 406894
rect 189822 406338 189854 406894
rect 189234 370894 189854 406338
rect 189234 370338 189266 370894
rect 189822 370338 189854 370894
rect 189234 334894 189854 370338
rect 189234 334338 189266 334894
rect 189822 334338 189854 334894
rect 189234 298894 189854 334338
rect 189234 298338 189266 298894
rect 189822 298338 189854 298894
rect 185168 270334 185488 270366
rect 185168 270098 185210 270334
rect 185446 270098 185488 270334
rect 185168 270014 185488 270098
rect 185168 269778 185210 270014
rect 185446 269778 185488 270014
rect 185168 269746 185488 269778
rect 181794 254898 181826 255454
rect 182382 254898 182414 255454
rect 177488 223174 177808 223206
rect 177488 222938 177530 223174
rect 177766 222938 177808 223174
rect 177488 222854 177808 222938
rect 177488 222618 177530 222854
rect 177766 222618 177808 222854
rect 177488 222586 177808 222618
rect 171834 208938 171866 209494
rect 172422 208938 172454 209494
rect 169808 183454 170128 183486
rect 169808 183218 169850 183454
rect 170086 183218 170128 183454
rect 169808 183134 170128 183218
rect 169808 182898 169850 183134
rect 170086 182898 170128 183134
rect 169808 182866 170128 182898
rect 168114 169218 168146 169774
rect 168702 169218 168734 169774
rect 168114 133774 168734 169218
rect 171834 173494 172454 208938
rect 181794 219454 182414 254898
rect 189234 262894 189854 298338
rect 192954 707718 193574 711590
rect 192954 707162 192986 707718
rect 193542 707162 193574 707718
rect 192954 698614 193574 707162
rect 192954 698058 192986 698614
rect 193542 698058 193574 698614
rect 192954 662614 193574 698058
rect 192954 662058 192986 662614
rect 193542 662058 193574 662614
rect 192954 626614 193574 662058
rect 192954 626058 192986 626614
rect 193542 626058 193574 626614
rect 192954 590614 193574 626058
rect 192954 590058 192986 590614
rect 193542 590058 193574 590614
rect 192954 554614 193574 590058
rect 192954 554058 192986 554614
rect 193542 554058 193574 554614
rect 192954 518614 193574 554058
rect 192954 518058 192986 518614
rect 193542 518058 193574 518614
rect 192954 482614 193574 518058
rect 192954 482058 192986 482614
rect 193542 482058 193574 482614
rect 192954 446614 193574 482058
rect 192954 446058 192986 446614
rect 193542 446058 193574 446614
rect 192954 410614 193574 446058
rect 192954 410058 192986 410614
rect 193542 410058 193574 410614
rect 192954 374614 193574 410058
rect 192954 374058 192986 374614
rect 193542 374058 193574 374614
rect 192954 338614 193574 374058
rect 192954 338058 192986 338614
rect 193542 338058 193574 338614
rect 192954 302614 193574 338058
rect 192954 302058 192986 302614
rect 193542 302058 193574 302614
rect 192954 282628 193574 302058
rect 196674 708678 197294 711590
rect 196674 708122 196706 708678
rect 197262 708122 197294 708678
rect 196674 666334 197294 708122
rect 196674 665778 196706 666334
rect 197262 665778 197294 666334
rect 196674 630334 197294 665778
rect 196674 629778 196706 630334
rect 197262 629778 197294 630334
rect 196674 594334 197294 629778
rect 196674 593778 196706 594334
rect 197262 593778 197294 594334
rect 196674 558334 197294 593778
rect 196674 557778 196706 558334
rect 197262 557778 197294 558334
rect 196674 522334 197294 557778
rect 196674 521778 196706 522334
rect 197262 521778 197294 522334
rect 196674 486334 197294 521778
rect 196674 485778 196706 486334
rect 197262 485778 197294 486334
rect 196674 450334 197294 485778
rect 196674 449778 196706 450334
rect 197262 449778 197294 450334
rect 196674 414334 197294 449778
rect 196674 413778 196706 414334
rect 197262 413778 197294 414334
rect 196674 378334 197294 413778
rect 196674 377778 196706 378334
rect 197262 377778 197294 378334
rect 196674 342334 197294 377778
rect 196674 341778 196706 342334
rect 197262 341778 197294 342334
rect 196674 306334 197294 341778
rect 196674 305778 196706 306334
rect 197262 305778 197294 306334
rect 192848 274054 193168 274086
rect 192848 273818 192890 274054
rect 193126 273818 193168 274054
rect 192848 273734 193168 273818
rect 192848 273498 192890 273734
rect 193126 273498 193168 273734
rect 192848 273466 193168 273498
rect 189234 262338 189266 262894
rect 189822 262338 189854 262894
rect 185168 234334 185488 234366
rect 185168 234098 185210 234334
rect 185446 234098 185488 234334
rect 185168 234014 185488 234098
rect 185168 233778 185210 234014
rect 185446 233778 185488 234014
rect 185168 233746 185488 233778
rect 181794 218898 181826 219454
rect 182382 218898 182414 219454
rect 177488 187174 177808 187206
rect 177488 186938 177530 187174
rect 177766 186938 177808 187174
rect 177488 186854 177808 186938
rect 177488 186618 177530 186854
rect 177766 186618 177808 186854
rect 177488 186586 177808 186618
rect 171834 172938 171866 173494
rect 172422 172938 172454 173494
rect 169808 147454 170128 147486
rect 169808 147218 169850 147454
rect 170086 147218 170128 147454
rect 169808 147134 170128 147218
rect 169808 146898 169850 147134
rect 170086 146898 170128 147134
rect 169808 146866 170128 146898
rect 168114 133218 168146 133774
rect 168702 133218 168734 133774
rect 168114 97774 168734 133218
rect 171834 137494 172454 172938
rect 181794 183454 182414 218898
rect 189234 226894 189854 262338
rect 196674 270334 197294 305778
rect 200394 709638 201014 711590
rect 200394 709082 200426 709638
rect 200982 709082 201014 709638
rect 200394 670054 201014 709082
rect 200394 669498 200426 670054
rect 200982 669498 201014 670054
rect 200394 634054 201014 669498
rect 200394 633498 200426 634054
rect 200982 633498 201014 634054
rect 200394 598054 201014 633498
rect 200394 597498 200426 598054
rect 200982 597498 201014 598054
rect 200394 562054 201014 597498
rect 200394 561498 200426 562054
rect 200982 561498 201014 562054
rect 200394 526054 201014 561498
rect 200394 525498 200426 526054
rect 200982 525498 201014 526054
rect 200394 490054 201014 525498
rect 200394 489498 200426 490054
rect 200982 489498 201014 490054
rect 200394 454054 201014 489498
rect 200394 453498 200426 454054
rect 200982 453498 201014 454054
rect 200394 418054 201014 453498
rect 200394 417498 200426 418054
rect 200982 417498 201014 418054
rect 200394 382054 201014 417498
rect 200394 381498 200426 382054
rect 200982 381498 201014 382054
rect 200394 346054 201014 381498
rect 200394 345498 200426 346054
rect 200982 345498 201014 346054
rect 200394 310054 201014 345498
rect 200394 309498 200426 310054
rect 200982 309498 201014 310054
rect 200394 282628 201014 309498
rect 204114 710598 204734 711590
rect 204114 710042 204146 710598
rect 204702 710042 204734 710598
rect 204114 673774 204734 710042
rect 204114 673218 204146 673774
rect 204702 673218 204734 673774
rect 204114 637774 204734 673218
rect 204114 637218 204146 637774
rect 204702 637218 204734 637774
rect 204114 601774 204734 637218
rect 204114 601218 204146 601774
rect 204702 601218 204734 601774
rect 204114 565774 204734 601218
rect 204114 565218 204146 565774
rect 204702 565218 204734 565774
rect 204114 529774 204734 565218
rect 204114 529218 204146 529774
rect 204702 529218 204734 529774
rect 204114 493774 204734 529218
rect 204114 493218 204146 493774
rect 204702 493218 204734 493774
rect 204114 457774 204734 493218
rect 204114 457218 204146 457774
rect 204702 457218 204734 457774
rect 204114 421774 204734 457218
rect 204114 421218 204146 421774
rect 204702 421218 204734 421774
rect 204114 385774 204734 421218
rect 204114 385218 204146 385774
rect 204702 385218 204734 385774
rect 204114 349774 204734 385218
rect 204114 349218 204146 349774
rect 204702 349218 204734 349774
rect 204114 313774 204734 349218
rect 204114 313218 204146 313774
rect 204702 313218 204734 313774
rect 196674 269778 196706 270334
rect 197262 269778 197294 270334
rect 192848 238054 193168 238086
rect 192848 237818 192890 238054
rect 193126 237818 193168 238054
rect 192848 237734 193168 237818
rect 192848 237498 192890 237734
rect 193126 237498 193168 237734
rect 192848 237466 193168 237498
rect 189234 226338 189266 226894
rect 189822 226338 189854 226894
rect 185168 198334 185488 198366
rect 185168 198098 185210 198334
rect 185446 198098 185488 198334
rect 185168 198014 185488 198098
rect 185168 197778 185210 198014
rect 185446 197778 185488 198014
rect 185168 197746 185488 197778
rect 181794 182898 181826 183454
rect 182382 182898 182414 183454
rect 177488 151174 177808 151206
rect 177488 150938 177530 151174
rect 177766 150938 177808 151174
rect 177488 150854 177808 150938
rect 177488 150618 177530 150854
rect 177766 150618 177808 150854
rect 177488 150586 177808 150618
rect 171834 136938 171866 137494
rect 172422 136938 172454 137494
rect 169808 111454 170128 111486
rect 169808 111218 169850 111454
rect 170086 111218 170128 111454
rect 169808 111134 170128 111218
rect 169808 110898 169850 111134
rect 170086 110898 170128 111134
rect 169808 110866 170128 110898
rect 168114 97218 168146 97774
rect 168702 97218 168734 97774
rect 168114 61774 168734 97218
rect 171834 101494 172454 136938
rect 181794 147454 182414 182898
rect 189234 190894 189854 226338
rect 196674 234334 197294 269778
rect 204114 277774 204734 313218
rect 207834 711558 208454 711590
rect 207834 711002 207866 711558
rect 208422 711002 208454 711558
rect 207834 677494 208454 711002
rect 207834 676938 207866 677494
rect 208422 676938 208454 677494
rect 207834 641494 208454 676938
rect 207834 640938 207866 641494
rect 208422 640938 208454 641494
rect 207834 605494 208454 640938
rect 207834 604938 207866 605494
rect 208422 604938 208454 605494
rect 207834 569494 208454 604938
rect 207834 568938 207866 569494
rect 208422 568938 208454 569494
rect 207834 533494 208454 568938
rect 207834 532938 207866 533494
rect 208422 532938 208454 533494
rect 207834 497494 208454 532938
rect 207834 496938 207866 497494
rect 208422 496938 208454 497494
rect 207834 461494 208454 496938
rect 207834 460938 207866 461494
rect 208422 460938 208454 461494
rect 207834 425494 208454 460938
rect 207834 424938 207866 425494
rect 208422 424938 208454 425494
rect 207834 389494 208454 424938
rect 207834 388938 207866 389494
rect 208422 388938 208454 389494
rect 207834 353494 208454 388938
rect 207834 352938 207866 353494
rect 208422 352938 208454 353494
rect 207834 317494 208454 352938
rect 207834 316938 207866 317494
rect 208422 316938 208454 317494
rect 207834 282628 208454 316938
rect 217794 704838 218414 711590
rect 217794 704282 217826 704838
rect 218382 704282 218414 704838
rect 217794 687454 218414 704282
rect 217794 686898 217826 687454
rect 218382 686898 218414 687454
rect 217794 651454 218414 686898
rect 217794 650898 217826 651454
rect 218382 650898 218414 651454
rect 217794 615454 218414 650898
rect 217794 614898 217826 615454
rect 218382 614898 218414 615454
rect 217794 579454 218414 614898
rect 217794 578898 217826 579454
rect 218382 578898 218414 579454
rect 217794 543454 218414 578898
rect 217794 542898 217826 543454
rect 218382 542898 218414 543454
rect 217794 507454 218414 542898
rect 217794 506898 217826 507454
rect 218382 506898 218414 507454
rect 217794 471454 218414 506898
rect 217794 470898 217826 471454
rect 218382 470898 218414 471454
rect 217794 435454 218414 470898
rect 217794 434898 217826 435454
rect 218382 434898 218414 435454
rect 217794 399454 218414 434898
rect 217794 398898 217826 399454
rect 218382 398898 218414 399454
rect 217794 363454 218414 398898
rect 217794 362898 217826 363454
rect 218382 362898 218414 363454
rect 217794 327454 218414 362898
rect 217794 326898 217826 327454
rect 218382 326898 218414 327454
rect 217794 291454 218414 326898
rect 217794 290898 217826 291454
rect 218382 290898 218414 291454
rect 204114 277218 204146 277774
rect 204702 277218 204734 277774
rect 200528 255454 200848 255486
rect 200528 255218 200570 255454
rect 200806 255218 200848 255454
rect 200528 255134 200848 255218
rect 200528 254898 200570 255134
rect 200806 254898 200848 255134
rect 200528 254866 200848 254898
rect 196674 233778 196706 234334
rect 197262 233778 197294 234334
rect 192848 202054 193168 202086
rect 192848 201818 192890 202054
rect 193126 201818 193168 202054
rect 192848 201734 193168 201818
rect 192848 201498 192890 201734
rect 193126 201498 193168 201734
rect 192848 201466 193168 201498
rect 189234 190338 189266 190894
rect 189822 190338 189854 190894
rect 185168 162334 185488 162366
rect 185168 162098 185210 162334
rect 185446 162098 185488 162334
rect 185168 162014 185488 162098
rect 185168 161778 185210 162014
rect 185446 161778 185488 162014
rect 185168 161746 185488 161778
rect 181794 146898 181826 147454
rect 182382 146898 182414 147454
rect 177488 115174 177808 115206
rect 177488 114938 177530 115174
rect 177766 114938 177808 115174
rect 177488 114854 177808 114938
rect 177488 114618 177530 114854
rect 177766 114618 177808 114854
rect 177488 114586 177808 114618
rect 171834 100938 171866 101494
rect 172422 100938 172454 101494
rect 169808 75454 170128 75486
rect 169808 75218 169850 75454
rect 170086 75218 170128 75454
rect 169808 75134 170128 75218
rect 169808 74898 169850 75134
rect 170086 74898 170128 75134
rect 169808 74866 170128 74898
rect 168114 61218 168146 61774
rect 168702 61218 168734 61774
rect 168114 25774 168734 61218
rect 171834 65494 172454 100938
rect 181794 111454 182414 146898
rect 189234 154894 189854 190338
rect 196674 198334 197294 233778
rect 204114 241774 204734 277218
rect 215888 270334 216208 270366
rect 215888 270098 215930 270334
rect 216166 270098 216208 270334
rect 215888 270014 216208 270098
rect 215888 269778 215930 270014
rect 216166 269778 216208 270014
rect 215888 269746 216208 269778
rect 208208 259174 208528 259206
rect 208208 258938 208250 259174
rect 208486 258938 208528 259174
rect 208208 258854 208528 258938
rect 208208 258618 208250 258854
rect 208486 258618 208528 258854
rect 208208 258586 208528 258618
rect 204114 241218 204146 241774
rect 204702 241218 204734 241774
rect 200528 219454 200848 219486
rect 200528 219218 200570 219454
rect 200806 219218 200848 219454
rect 200528 219134 200848 219218
rect 200528 218898 200570 219134
rect 200806 218898 200848 219134
rect 200528 218866 200848 218898
rect 196674 197778 196706 198334
rect 197262 197778 197294 198334
rect 192848 166054 193168 166086
rect 192848 165818 192890 166054
rect 193126 165818 193168 166054
rect 192848 165734 193168 165818
rect 192848 165498 192890 165734
rect 193126 165498 193168 165734
rect 192848 165466 193168 165498
rect 189234 154338 189266 154894
rect 189822 154338 189854 154894
rect 185168 126334 185488 126366
rect 185168 126098 185210 126334
rect 185446 126098 185488 126334
rect 185168 126014 185488 126098
rect 185168 125778 185210 126014
rect 185446 125778 185488 126014
rect 185168 125746 185488 125778
rect 181794 110898 181826 111454
rect 182382 110898 182414 111454
rect 177488 79174 177808 79206
rect 177488 78938 177530 79174
rect 177766 78938 177808 79174
rect 177488 78854 177808 78938
rect 177488 78618 177530 78854
rect 177766 78618 177808 78854
rect 177488 78586 177808 78618
rect 171834 64938 171866 65494
rect 172422 64938 172454 65494
rect 169808 39454 170128 39486
rect 169808 39218 169850 39454
rect 170086 39218 170128 39454
rect 169808 39134 170128 39218
rect 169808 38898 169850 39134
rect 170086 38898 170128 39134
rect 169808 38866 170128 38898
rect 168114 25218 168146 25774
rect 168702 25218 168734 25774
rect 168114 -6106 168734 25218
rect 168114 -6662 168146 -6106
rect 168702 -6662 168734 -6106
rect 168114 -7654 168734 -6662
rect 171834 29494 172454 64938
rect 181794 75454 182414 110898
rect 189234 118894 189854 154338
rect 196674 162334 197294 197778
rect 204114 205774 204734 241218
rect 217794 255454 218414 290898
rect 217794 254898 217826 255454
rect 218382 254898 218414 255454
rect 215888 234334 216208 234366
rect 215888 234098 215930 234334
rect 216166 234098 216208 234334
rect 215888 234014 216208 234098
rect 215888 233778 215930 234014
rect 216166 233778 216208 234014
rect 215888 233746 216208 233778
rect 208208 223174 208528 223206
rect 208208 222938 208250 223174
rect 208486 222938 208528 223174
rect 208208 222854 208528 222938
rect 208208 222618 208250 222854
rect 208486 222618 208528 222854
rect 208208 222586 208528 222618
rect 204114 205218 204146 205774
rect 204702 205218 204734 205774
rect 200528 183454 200848 183486
rect 200528 183218 200570 183454
rect 200806 183218 200848 183454
rect 200528 183134 200848 183218
rect 200528 182898 200570 183134
rect 200806 182898 200848 183134
rect 200528 182866 200848 182898
rect 196674 161778 196706 162334
rect 197262 161778 197294 162334
rect 192848 130054 193168 130086
rect 192848 129818 192890 130054
rect 193126 129818 193168 130054
rect 192848 129734 193168 129818
rect 192848 129498 192890 129734
rect 193126 129498 193168 129734
rect 192848 129466 193168 129498
rect 189234 118338 189266 118894
rect 189822 118338 189854 118894
rect 185168 90334 185488 90366
rect 185168 90098 185210 90334
rect 185446 90098 185488 90334
rect 185168 90014 185488 90098
rect 185168 89778 185210 90014
rect 185446 89778 185488 90014
rect 185168 89746 185488 89778
rect 181794 74898 181826 75454
rect 182382 74898 182414 75454
rect 177488 43174 177808 43206
rect 177488 42938 177530 43174
rect 177766 42938 177808 43174
rect 177488 42854 177808 42938
rect 177488 42618 177530 42854
rect 177766 42618 177808 42854
rect 177488 42586 177808 42618
rect 171834 28938 171866 29494
rect 172422 28938 172454 29494
rect 171834 -7066 172454 28938
rect 181794 39454 182414 74898
rect 189234 82894 189854 118338
rect 196674 126334 197294 161778
rect 204114 169774 204734 205218
rect 217794 219454 218414 254898
rect 217794 218898 217826 219454
rect 218382 218898 218414 219454
rect 215888 198334 216208 198366
rect 215888 198098 215930 198334
rect 216166 198098 216208 198334
rect 215888 198014 216208 198098
rect 215888 197778 215930 198014
rect 216166 197778 216208 198014
rect 215888 197746 216208 197778
rect 208208 187174 208528 187206
rect 208208 186938 208250 187174
rect 208486 186938 208528 187174
rect 208208 186854 208528 186938
rect 208208 186618 208250 186854
rect 208486 186618 208528 186854
rect 208208 186586 208528 186618
rect 204114 169218 204146 169774
rect 204702 169218 204734 169774
rect 200528 147454 200848 147486
rect 200528 147218 200570 147454
rect 200806 147218 200848 147454
rect 200528 147134 200848 147218
rect 200528 146898 200570 147134
rect 200806 146898 200848 147134
rect 200528 146866 200848 146898
rect 196674 125778 196706 126334
rect 197262 125778 197294 126334
rect 192848 94054 193168 94086
rect 192848 93818 192890 94054
rect 193126 93818 193168 94054
rect 192848 93734 193168 93818
rect 192848 93498 192890 93734
rect 193126 93498 193168 93734
rect 192848 93466 193168 93498
rect 189234 82338 189266 82894
rect 189822 82338 189854 82894
rect 185168 54334 185488 54366
rect 185168 54098 185210 54334
rect 185446 54098 185488 54334
rect 185168 54014 185488 54098
rect 185168 53778 185210 54014
rect 185446 53778 185488 54014
rect 185168 53746 185488 53778
rect 181794 38898 181826 39454
rect 182382 38898 182414 39454
rect 177488 7174 177808 7206
rect 177488 6938 177530 7174
rect 177766 6938 177808 7174
rect 177488 6854 177808 6938
rect 177488 6618 177530 6854
rect 177766 6618 177808 6854
rect 177488 6586 177808 6618
rect 171834 -7622 171866 -7066
rect 172422 -7622 172454 -7066
rect 171834 -7654 172454 -7622
rect 181794 3454 182414 38898
rect 189234 46894 189854 82338
rect 196674 90334 197294 125778
rect 204114 133774 204734 169218
rect 217794 183454 218414 218898
rect 217794 182898 217826 183454
rect 218382 182898 218414 183454
rect 215888 162334 216208 162366
rect 215888 162098 215930 162334
rect 216166 162098 216208 162334
rect 215888 162014 216208 162098
rect 215888 161778 215930 162014
rect 216166 161778 216208 162014
rect 215888 161746 216208 161778
rect 208208 151174 208528 151206
rect 208208 150938 208250 151174
rect 208486 150938 208528 151174
rect 208208 150854 208528 150938
rect 208208 150618 208250 150854
rect 208486 150618 208528 150854
rect 208208 150586 208528 150618
rect 204114 133218 204146 133774
rect 204702 133218 204734 133774
rect 200528 111454 200848 111486
rect 200528 111218 200570 111454
rect 200806 111218 200848 111454
rect 200528 111134 200848 111218
rect 200528 110898 200570 111134
rect 200806 110898 200848 111134
rect 200528 110866 200848 110898
rect 196674 89778 196706 90334
rect 197262 89778 197294 90334
rect 192848 58054 193168 58086
rect 192848 57818 192890 58054
rect 193126 57818 193168 58054
rect 192848 57734 193168 57818
rect 192848 57498 192890 57734
rect 193126 57498 193168 57734
rect 192848 57466 193168 57498
rect 189234 46338 189266 46894
rect 189822 46338 189854 46894
rect 185168 18334 185488 18366
rect 185168 18098 185210 18334
rect 185446 18098 185488 18334
rect 185168 18014 185488 18098
rect 185168 17778 185210 18014
rect 185446 17778 185488 18014
rect 185168 17746 185488 17778
rect 181794 2898 181826 3454
rect 182382 2898 182414 3454
rect 189234 10894 189854 46338
rect 196674 54334 197294 89778
rect 204114 97774 204734 133218
rect 217794 147454 218414 182898
rect 217794 146898 217826 147454
rect 218382 146898 218414 147454
rect 215888 126334 216208 126366
rect 215888 126098 215930 126334
rect 216166 126098 216208 126334
rect 215888 126014 216208 126098
rect 215888 125778 215930 126014
rect 216166 125778 216208 126014
rect 215888 125746 216208 125778
rect 208208 115174 208528 115206
rect 208208 114938 208250 115174
rect 208486 114938 208528 115174
rect 208208 114854 208528 114938
rect 208208 114618 208250 114854
rect 208486 114618 208528 114854
rect 208208 114586 208528 114618
rect 204114 97218 204146 97774
rect 204702 97218 204734 97774
rect 200528 75454 200848 75486
rect 200528 75218 200570 75454
rect 200806 75218 200848 75454
rect 200528 75134 200848 75218
rect 200528 74898 200570 75134
rect 200806 74898 200848 75134
rect 200528 74866 200848 74898
rect 196674 53778 196706 54334
rect 197262 53778 197294 54334
rect 192848 22054 193168 22086
rect 192848 21818 192890 22054
rect 193126 21818 193168 22054
rect 192848 21734 193168 21818
rect 192848 21498 192890 21734
rect 193126 21498 193168 21734
rect 192848 21466 193168 21498
rect 189234 10338 189266 10894
rect 189822 10338 189854 10894
rect 181794 -346 182414 2898
rect 181794 -902 181826 -346
rect 182382 -902 182414 -346
rect 181794 -7654 182414 -902
rect 185514 -1306 186134 2988
rect 185514 -1862 185546 -1306
rect 186102 -1862 186134 -1306
rect 185514 -7654 186134 -1862
rect 189234 -2266 189854 10338
rect 196674 18334 197294 53778
rect 204114 61774 204734 97218
rect 217794 111454 218414 146898
rect 217794 110898 217826 111454
rect 218382 110898 218414 111454
rect 215888 90334 216208 90366
rect 215888 90098 215930 90334
rect 216166 90098 216208 90334
rect 215888 90014 216208 90098
rect 215888 89778 215930 90014
rect 216166 89778 216208 90014
rect 215888 89746 216208 89778
rect 208208 79174 208528 79206
rect 208208 78938 208250 79174
rect 208486 78938 208528 79174
rect 208208 78854 208528 78938
rect 208208 78618 208250 78854
rect 208486 78618 208528 78854
rect 208208 78586 208528 78618
rect 204114 61218 204146 61774
rect 204702 61218 204734 61774
rect 200528 39454 200848 39486
rect 200528 39218 200570 39454
rect 200806 39218 200848 39454
rect 200528 39134 200848 39218
rect 200528 38898 200570 39134
rect 200806 38898 200848 39134
rect 200528 38866 200848 38898
rect 196674 17778 196706 18334
rect 197262 17778 197294 18334
rect 189234 -2822 189266 -2266
rect 189822 -2822 189854 -2266
rect 189234 -7654 189854 -2822
rect 192954 -3226 193574 2988
rect 192954 -3782 192986 -3226
rect 193542 -3782 193574 -3226
rect 192954 -7654 193574 -3782
rect 196674 -4186 197294 17778
rect 204114 25774 204734 61218
rect 217794 75454 218414 110898
rect 217794 74898 217826 75454
rect 218382 74898 218414 75454
rect 215888 54334 216208 54366
rect 215888 54098 215930 54334
rect 216166 54098 216208 54334
rect 215888 54014 216208 54098
rect 215888 53778 215930 54014
rect 216166 53778 216208 54014
rect 215888 53746 216208 53778
rect 208208 43174 208528 43206
rect 208208 42938 208250 43174
rect 208486 42938 208528 43174
rect 208208 42854 208528 42938
rect 208208 42618 208250 42854
rect 208486 42618 208528 42854
rect 208208 42586 208528 42618
rect 204114 25218 204146 25774
rect 204702 25218 204734 25774
rect 196674 -4742 196706 -4186
rect 197262 -4742 197294 -4186
rect 196674 -7654 197294 -4742
rect 200394 -5146 201014 2988
rect 200394 -5702 200426 -5146
rect 200982 -5702 201014 -5146
rect 200394 -7654 201014 -5702
rect 204114 -6106 204734 25218
rect 217794 39454 218414 74898
rect 217794 38898 217826 39454
rect 218382 38898 218414 39454
rect 215888 18334 216208 18366
rect 215888 18098 215930 18334
rect 216166 18098 216208 18334
rect 215888 18014 216208 18098
rect 215888 17778 215930 18014
rect 216166 17778 216208 18014
rect 215888 17746 216208 17778
rect 208208 7174 208528 7206
rect 208208 6938 208250 7174
rect 208486 6938 208528 7174
rect 208208 6854 208528 6938
rect 208208 6618 208250 6854
rect 208486 6618 208528 6854
rect 208208 6586 208528 6618
rect 217794 3454 218414 38898
rect 204114 -6662 204146 -6106
rect 204702 -6662 204734 -6106
rect 204114 -7654 204734 -6662
rect 207834 -7066 208454 2988
rect 207834 -7622 207866 -7066
rect 208422 -7622 208454 -7066
rect 207834 -7654 208454 -7622
rect 217794 2898 217826 3454
rect 218382 2898 218414 3454
rect 217794 -346 218414 2898
rect 217794 -902 217826 -346
rect 218382 -902 218414 -346
rect 217794 -7654 218414 -902
rect 221514 705798 222134 711590
rect 221514 705242 221546 705798
rect 222102 705242 222134 705798
rect 221514 691174 222134 705242
rect 221514 690618 221546 691174
rect 222102 690618 222134 691174
rect 221514 655174 222134 690618
rect 221514 654618 221546 655174
rect 222102 654618 222134 655174
rect 221514 619174 222134 654618
rect 221514 618618 221546 619174
rect 222102 618618 222134 619174
rect 221514 583174 222134 618618
rect 221514 582618 221546 583174
rect 222102 582618 222134 583174
rect 221514 547174 222134 582618
rect 221514 546618 221546 547174
rect 222102 546618 222134 547174
rect 221514 511174 222134 546618
rect 221514 510618 221546 511174
rect 222102 510618 222134 511174
rect 221514 475174 222134 510618
rect 221514 474618 221546 475174
rect 222102 474618 222134 475174
rect 221514 439174 222134 474618
rect 221514 438618 221546 439174
rect 222102 438618 222134 439174
rect 221514 403174 222134 438618
rect 221514 402618 221546 403174
rect 222102 402618 222134 403174
rect 221514 367174 222134 402618
rect 221514 366618 221546 367174
rect 222102 366618 222134 367174
rect 221514 331174 222134 366618
rect 221514 330618 221546 331174
rect 222102 330618 222134 331174
rect 221514 295174 222134 330618
rect 221514 294618 221546 295174
rect 222102 294618 222134 295174
rect 221514 259174 222134 294618
rect 225234 706758 225854 711590
rect 225234 706202 225266 706758
rect 225822 706202 225854 706758
rect 225234 694894 225854 706202
rect 225234 694338 225266 694894
rect 225822 694338 225854 694894
rect 225234 658894 225854 694338
rect 225234 658338 225266 658894
rect 225822 658338 225854 658894
rect 225234 622894 225854 658338
rect 225234 622338 225266 622894
rect 225822 622338 225854 622894
rect 225234 586894 225854 622338
rect 225234 586338 225266 586894
rect 225822 586338 225854 586894
rect 225234 550894 225854 586338
rect 225234 550338 225266 550894
rect 225822 550338 225854 550894
rect 225234 514894 225854 550338
rect 225234 514338 225266 514894
rect 225822 514338 225854 514894
rect 225234 478894 225854 514338
rect 225234 478338 225266 478894
rect 225822 478338 225854 478894
rect 225234 442894 225854 478338
rect 225234 442338 225266 442894
rect 225822 442338 225854 442894
rect 225234 406894 225854 442338
rect 225234 406338 225266 406894
rect 225822 406338 225854 406894
rect 225234 370894 225854 406338
rect 225234 370338 225266 370894
rect 225822 370338 225854 370894
rect 225234 334894 225854 370338
rect 225234 334338 225266 334894
rect 225822 334338 225854 334894
rect 225234 298894 225854 334338
rect 225234 298338 225266 298894
rect 225822 298338 225854 298894
rect 223568 274054 223888 274086
rect 223568 273818 223610 274054
rect 223846 273818 223888 274054
rect 223568 273734 223888 273818
rect 223568 273498 223610 273734
rect 223846 273498 223888 273734
rect 223568 273466 223888 273498
rect 221514 258618 221546 259174
rect 222102 258618 222134 259174
rect 221514 223174 222134 258618
rect 225234 262894 225854 298338
rect 225234 262338 225266 262894
rect 225822 262338 225854 262894
rect 223568 238054 223888 238086
rect 223568 237818 223610 238054
rect 223846 237818 223888 238054
rect 223568 237734 223888 237818
rect 223568 237498 223610 237734
rect 223846 237498 223888 237734
rect 223568 237466 223888 237498
rect 221514 222618 221546 223174
rect 222102 222618 222134 223174
rect 221514 187174 222134 222618
rect 225234 226894 225854 262338
rect 225234 226338 225266 226894
rect 225822 226338 225854 226894
rect 223568 202054 223888 202086
rect 223568 201818 223610 202054
rect 223846 201818 223888 202054
rect 223568 201734 223888 201818
rect 223568 201498 223610 201734
rect 223846 201498 223888 201734
rect 223568 201466 223888 201498
rect 221514 186618 221546 187174
rect 222102 186618 222134 187174
rect 221514 151174 222134 186618
rect 225234 190894 225854 226338
rect 225234 190338 225266 190894
rect 225822 190338 225854 190894
rect 223568 166054 223888 166086
rect 223568 165818 223610 166054
rect 223846 165818 223888 166054
rect 223568 165734 223888 165818
rect 223568 165498 223610 165734
rect 223846 165498 223888 165734
rect 223568 165466 223888 165498
rect 221514 150618 221546 151174
rect 222102 150618 222134 151174
rect 221514 115174 222134 150618
rect 225234 154894 225854 190338
rect 225234 154338 225266 154894
rect 225822 154338 225854 154894
rect 223568 130054 223888 130086
rect 223568 129818 223610 130054
rect 223846 129818 223888 130054
rect 223568 129734 223888 129818
rect 223568 129498 223610 129734
rect 223846 129498 223888 129734
rect 223568 129466 223888 129498
rect 221514 114618 221546 115174
rect 222102 114618 222134 115174
rect 221514 79174 222134 114618
rect 225234 118894 225854 154338
rect 225234 118338 225266 118894
rect 225822 118338 225854 118894
rect 223568 94054 223888 94086
rect 223568 93818 223610 94054
rect 223846 93818 223888 94054
rect 223568 93734 223888 93818
rect 223568 93498 223610 93734
rect 223846 93498 223888 93734
rect 223568 93466 223888 93498
rect 221514 78618 221546 79174
rect 222102 78618 222134 79174
rect 221514 43174 222134 78618
rect 225234 82894 225854 118338
rect 225234 82338 225266 82894
rect 225822 82338 225854 82894
rect 223568 58054 223888 58086
rect 223568 57818 223610 58054
rect 223846 57818 223888 58054
rect 223568 57734 223888 57818
rect 223568 57498 223610 57734
rect 223846 57498 223888 57734
rect 223568 57466 223888 57498
rect 221514 42618 221546 43174
rect 222102 42618 222134 43174
rect 221514 7174 222134 42618
rect 225234 46894 225854 82338
rect 225234 46338 225266 46894
rect 225822 46338 225854 46894
rect 223568 22054 223888 22086
rect 223568 21818 223610 22054
rect 223846 21818 223888 22054
rect 223568 21734 223888 21818
rect 223568 21498 223610 21734
rect 223846 21498 223888 21734
rect 223568 21466 223888 21498
rect 221514 6618 221546 7174
rect 222102 6618 222134 7174
rect 221514 -1306 222134 6618
rect 221514 -1862 221546 -1306
rect 222102 -1862 222134 -1306
rect 221514 -7654 222134 -1862
rect 225234 10894 225854 46338
rect 225234 10338 225266 10894
rect 225822 10338 225854 10894
rect 225234 -2266 225854 10338
rect 225234 -2822 225266 -2266
rect 225822 -2822 225854 -2266
rect 225234 -7654 225854 -2822
rect 228954 707718 229574 711590
rect 228954 707162 228986 707718
rect 229542 707162 229574 707718
rect 228954 698614 229574 707162
rect 228954 698058 228986 698614
rect 229542 698058 229574 698614
rect 228954 662614 229574 698058
rect 228954 662058 228986 662614
rect 229542 662058 229574 662614
rect 228954 626614 229574 662058
rect 228954 626058 228986 626614
rect 229542 626058 229574 626614
rect 228954 590614 229574 626058
rect 228954 590058 228986 590614
rect 229542 590058 229574 590614
rect 228954 554614 229574 590058
rect 228954 554058 228986 554614
rect 229542 554058 229574 554614
rect 228954 518614 229574 554058
rect 228954 518058 228986 518614
rect 229542 518058 229574 518614
rect 228954 482614 229574 518058
rect 228954 482058 228986 482614
rect 229542 482058 229574 482614
rect 228954 446614 229574 482058
rect 228954 446058 228986 446614
rect 229542 446058 229574 446614
rect 228954 410614 229574 446058
rect 228954 410058 228986 410614
rect 229542 410058 229574 410614
rect 228954 374614 229574 410058
rect 228954 374058 228986 374614
rect 229542 374058 229574 374614
rect 228954 338614 229574 374058
rect 228954 338058 228986 338614
rect 229542 338058 229574 338614
rect 228954 302614 229574 338058
rect 228954 302058 228986 302614
rect 229542 302058 229574 302614
rect 228954 266614 229574 302058
rect 228954 266058 228986 266614
rect 229542 266058 229574 266614
rect 228954 230614 229574 266058
rect 232674 708678 233294 711590
rect 232674 708122 232706 708678
rect 233262 708122 233294 708678
rect 232674 666334 233294 708122
rect 232674 665778 232706 666334
rect 233262 665778 233294 666334
rect 232674 630334 233294 665778
rect 232674 629778 232706 630334
rect 233262 629778 233294 630334
rect 232674 594334 233294 629778
rect 232674 593778 232706 594334
rect 233262 593778 233294 594334
rect 232674 558334 233294 593778
rect 232674 557778 232706 558334
rect 233262 557778 233294 558334
rect 232674 522334 233294 557778
rect 232674 521778 232706 522334
rect 233262 521778 233294 522334
rect 232674 486334 233294 521778
rect 232674 485778 232706 486334
rect 233262 485778 233294 486334
rect 232674 450334 233294 485778
rect 232674 449778 232706 450334
rect 233262 449778 233294 450334
rect 232674 414334 233294 449778
rect 232674 413778 232706 414334
rect 233262 413778 233294 414334
rect 232674 378334 233294 413778
rect 232674 377778 232706 378334
rect 233262 377778 233294 378334
rect 232674 342334 233294 377778
rect 232674 341778 232706 342334
rect 233262 341778 233294 342334
rect 232674 306334 233294 341778
rect 232674 305778 232706 306334
rect 233262 305778 233294 306334
rect 232674 270334 233294 305778
rect 232674 269778 232706 270334
rect 233262 269778 233294 270334
rect 231248 255454 231568 255486
rect 231248 255218 231290 255454
rect 231526 255218 231568 255454
rect 231248 255134 231568 255218
rect 231248 254898 231290 255134
rect 231526 254898 231568 255134
rect 231248 254866 231568 254898
rect 228954 230058 228986 230614
rect 229542 230058 229574 230614
rect 228954 194614 229574 230058
rect 232674 234334 233294 269778
rect 232674 233778 232706 234334
rect 233262 233778 233294 234334
rect 231248 219454 231568 219486
rect 231248 219218 231290 219454
rect 231526 219218 231568 219454
rect 231248 219134 231568 219218
rect 231248 218898 231290 219134
rect 231526 218898 231568 219134
rect 231248 218866 231568 218898
rect 228954 194058 228986 194614
rect 229542 194058 229574 194614
rect 228954 158614 229574 194058
rect 232674 198334 233294 233778
rect 232674 197778 232706 198334
rect 233262 197778 233294 198334
rect 231248 183454 231568 183486
rect 231248 183218 231290 183454
rect 231526 183218 231568 183454
rect 231248 183134 231568 183218
rect 231248 182898 231290 183134
rect 231526 182898 231568 183134
rect 231248 182866 231568 182898
rect 228954 158058 228986 158614
rect 229542 158058 229574 158614
rect 228954 122614 229574 158058
rect 232674 162334 233294 197778
rect 232674 161778 232706 162334
rect 233262 161778 233294 162334
rect 231248 147454 231568 147486
rect 231248 147218 231290 147454
rect 231526 147218 231568 147454
rect 231248 147134 231568 147218
rect 231248 146898 231290 147134
rect 231526 146898 231568 147134
rect 231248 146866 231568 146898
rect 228954 122058 228986 122614
rect 229542 122058 229574 122614
rect 228954 86614 229574 122058
rect 232674 126334 233294 161778
rect 232674 125778 232706 126334
rect 233262 125778 233294 126334
rect 231248 111454 231568 111486
rect 231248 111218 231290 111454
rect 231526 111218 231568 111454
rect 231248 111134 231568 111218
rect 231248 110898 231290 111134
rect 231526 110898 231568 111134
rect 231248 110866 231568 110898
rect 228954 86058 228986 86614
rect 229542 86058 229574 86614
rect 228954 50614 229574 86058
rect 232674 90334 233294 125778
rect 232674 89778 232706 90334
rect 233262 89778 233294 90334
rect 231248 75454 231568 75486
rect 231248 75218 231290 75454
rect 231526 75218 231568 75454
rect 231248 75134 231568 75218
rect 231248 74898 231290 75134
rect 231526 74898 231568 75134
rect 231248 74866 231568 74898
rect 228954 50058 228986 50614
rect 229542 50058 229574 50614
rect 228954 14614 229574 50058
rect 232674 54334 233294 89778
rect 232674 53778 232706 54334
rect 233262 53778 233294 54334
rect 231248 39454 231568 39486
rect 231248 39218 231290 39454
rect 231526 39218 231568 39454
rect 231248 39134 231568 39218
rect 231248 38898 231290 39134
rect 231526 38898 231568 39134
rect 231248 38866 231568 38898
rect 228954 14058 228986 14614
rect 229542 14058 229574 14614
rect 228954 -3226 229574 14058
rect 228954 -3782 228986 -3226
rect 229542 -3782 229574 -3226
rect 228954 -7654 229574 -3782
rect 232674 18334 233294 53778
rect 232674 17778 232706 18334
rect 233262 17778 233294 18334
rect 232674 -4186 233294 17778
rect 232674 -4742 232706 -4186
rect 233262 -4742 233294 -4186
rect 232674 -7654 233294 -4742
rect 236394 709638 237014 711590
rect 236394 709082 236426 709638
rect 236982 709082 237014 709638
rect 236394 670054 237014 709082
rect 236394 669498 236426 670054
rect 236982 669498 237014 670054
rect 236394 634054 237014 669498
rect 236394 633498 236426 634054
rect 236982 633498 237014 634054
rect 236394 598054 237014 633498
rect 236394 597498 236426 598054
rect 236982 597498 237014 598054
rect 236394 562054 237014 597498
rect 236394 561498 236426 562054
rect 236982 561498 237014 562054
rect 236394 526054 237014 561498
rect 236394 525498 236426 526054
rect 236982 525498 237014 526054
rect 236394 490054 237014 525498
rect 236394 489498 236426 490054
rect 236982 489498 237014 490054
rect 236394 454054 237014 489498
rect 236394 453498 236426 454054
rect 236982 453498 237014 454054
rect 236394 418054 237014 453498
rect 236394 417498 236426 418054
rect 236982 417498 237014 418054
rect 236394 382054 237014 417498
rect 236394 381498 236426 382054
rect 236982 381498 237014 382054
rect 236394 346054 237014 381498
rect 236394 345498 236426 346054
rect 236982 345498 237014 346054
rect 236394 310054 237014 345498
rect 236394 309498 236426 310054
rect 236982 309498 237014 310054
rect 236394 274054 237014 309498
rect 236394 273498 236426 274054
rect 236982 273498 237014 274054
rect 236394 238054 237014 273498
rect 240114 710598 240734 711590
rect 240114 710042 240146 710598
rect 240702 710042 240734 710598
rect 240114 673774 240734 710042
rect 240114 673218 240146 673774
rect 240702 673218 240734 673774
rect 240114 637774 240734 673218
rect 240114 637218 240146 637774
rect 240702 637218 240734 637774
rect 240114 601774 240734 637218
rect 240114 601218 240146 601774
rect 240702 601218 240734 601774
rect 240114 565774 240734 601218
rect 240114 565218 240146 565774
rect 240702 565218 240734 565774
rect 240114 529774 240734 565218
rect 240114 529218 240146 529774
rect 240702 529218 240734 529774
rect 240114 493774 240734 529218
rect 240114 493218 240146 493774
rect 240702 493218 240734 493774
rect 240114 457774 240734 493218
rect 240114 457218 240146 457774
rect 240702 457218 240734 457774
rect 240114 421774 240734 457218
rect 240114 421218 240146 421774
rect 240702 421218 240734 421774
rect 240114 385774 240734 421218
rect 240114 385218 240146 385774
rect 240702 385218 240734 385774
rect 240114 349774 240734 385218
rect 240114 349218 240146 349774
rect 240702 349218 240734 349774
rect 240114 313774 240734 349218
rect 240114 313218 240146 313774
rect 240702 313218 240734 313774
rect 240114 277774 240734 313218
rect 240114 277218 240146 277774
rect 240702 277218 240734 277774
rect 238928 259174 239248 259206
rect 238928 258938 238970 259174
rect 239206 258938 239248 259174
rect 238928 258854 239248 258938
rect 238928 258618 238970 258854
rect 239206 258618 239248 258854
rect 238928 258586 239248 258618
rect 236394 237498 236426 238054
rect 236982 237498 237014 238054
rect 236394 202054 237014 237498
rect 240114 241774 240734 277218
rect 240114 241218 240146 241774
rect 240702 241218 240734 241774
rect 238928 223174 239248 223206
rect 238928 222938 238970 223174
rect 239206 222938 239248 223174
rect 238928 222854 239248 222938
rect 238928 222618 238970 222854
rect 239206 222618 239248 222854
rect 238928 222586 239248 222618
rect 236394 201498 236426 202054
rect 236982 201498 237014 202054
rect 236394 166054 237014 201498
rect 240114 205774 240734 241218
rect 240114 205218 240146 205774
rect 240702 205218 240734 205774
rect 238928 187174 239248 187206
rect 238928 186938 238970 187174
rect 239206 186938 239248 187174
rect 238928 186854 239248 186938
rect 238928 186618 238970 186854
rect 239206 186618 239248 186854
rect 238928 186586 239248 186618
rect 236394 165498 236426 166054
rect 236982 165498 237014 166054
rect 236394 130054 237014 165498
rect 240114 169774 240734 205218
rect 240114 169218 240146 169774
rect 240702 169218 240734 169774
rect 238928 151174 239248 151206
rect 238928 150938 238970 151174
rect 239206 150938 239248 151174
rect 238928 150854 239248 150938
rect 238928 150618 238970 150854
rect 239206 150618 239248 150854
rect 238928 150586 239248 150618
rect 236394 129498 236426 130054
rect 236982 129498 237014 130054
rect 236394 94054 237014 129498
rect 240114 133774 240734 169218
rect 240114 133218 240146 133774
rect 240702 133218 240734 133774
rect 238928 115174 239248 115206
rect 238928 114938 238970 115174
rect 239206 114938 239248 115174
rect 238928 114854 239248 114938
rect 238928 114618 238970 114854
rect 239206 114618 239248 114854
rect 238928 114586 239248 114618
rect 236394 93498 236426 94054
rect 236982 93498 237014 94054
rect 236394 58054 237014 93498
rect 240114 97774 240734 133218
rect 240114 97218 240146 97774
rect 240702 97218 240734 97774
rect 238928 79174 239248 79206
rect 238928 78938 238970 79174
rect 239206 78938 239248 79174
rect 238928 78854 239248 78938
rect 238928 78618 238970 78854
rect 239206 78618 239248 78854
rect 238928 78586 239248 78618
rect 236394 57498 236426 58054
rect 236982 57498 237014 58054
rect 236394 22054 237014 57498
rect 240114 61774 240734 97218
rect 240114 61218 240146 61774
rect 240702 61218 240734 61774
rect 238928 43174 239248 43206
rect 238928 42938 238970 43174
rect 239206 42938 239248 43174
rect 238928 42854 239248 42938
rect 238928 42618 238970 42854
rect 239206 42618 239248 42854
rect 238928 42586 239248 42618
rect 236394 21498 236426 22054
rect 236982 21498 237014 22054
rect 236394 -5146 237014 21498
rect 240114 25774 240734 61218
rect 240114 25218 240146 25774
rect 240702 25218 240734 25774
rect 238928 7174 239248 7206
rect 238928 6938 238970 7174
rect 239206 6938 239248 7174
rect 238928 6854 239248 6938
rect 238928 6618 238970 6854
rect 239206 6618 239248 6854
rect 238928 6586 239248 6618
rect 236394 -5702 236426 -5146
rect 236982 -5702 237014 -5146
rect 236394 -7654 237014 -5702
rect 240114 -6106 240734 25218
rect 240114 -6662 240146 -6106
rect 240702 -6662 240734 -6106
rect 240114 -7654 240734 -6662
rect 243834 711558 244454 711590
rect 243834 711002 243866 711558
rect 244422 711002 244454 711558
rect 243834 677494 244454 711002
rect 243834 676938 243866 677494
rect 244422 676938 244454 677494
rect 243834 641494 244454 676938
rect 243834 640938 243866 641494
rect 244422 640938 244454 641494
rect 243834 605494 244454 640938
rect 243834 604938 243866 605494
rect 244422 604938 244454 605494
rect 243834 569494 244454 604938
rect 243834 568938 243866 569494
rect 244422 568938 244454 569494
rect 243834 533494 244454 568938
rect 243834 532938 243866 533494
rect 244422 532938 244454 533494
rect 243834 497494 244454 532938
rect 243834 496938 243866 497494
rect 244422 496938 244454 497494
rect 243834 461494 244454 496938
rect 243834 460938 243866 461494
rect 244422 460938 244454 461494
rect 243834 425494 244454 460938
rect 243834 424938 243866 425494
rect 244422 424938 244454 425494
rect 243834 389494 244454 424938
rect 243834 388938 243866 389494
rect 244422 388938 244454 389494
rect 243834 353494 244454 388938
rect 243834 352938 243866 353494
rect 244422 352938 244454 353494
rect 243834 317494 244454 352938
rect 243834 316938 243866 317494
rect 244422 316938 244454 317494
rect 243834 281494 244454 316938
rect 253794 704838 254414 711590
rect 253794 704282 253826 704838
rect 254382 704282 254414 704838
rect 253794 687454 254414 704282
rect 253794 686898 253826 687454
rect 254382 686898 254414 687454
rect 253794 651454 254414 686898
rect 253794 650898 253826 651454
rect 254382 650898 254414 651454
rect 253794 615454 254414 650898
rect 253794 614898 253826 615454
rect 254382 614898 254414 615454
rect 253794 579454 254414 614898
rect 253794 578898 253826 579454
rect 254382 578898 254414 579454
rect 253794 543454 254414 578898
rect 253794 542898 253826 543454
rect 254382 542898 254414 543454
rect 253794 507454 254414 542898
rect 253794 506898 253826 507454
rect 254382 506898 254414 507454
rect 253794 471454 254414 506898
rect 253794 470898 253826 471454
rect 254382 470898 254414 471454
rect 253794 435454 254414 470898
rect 253794 434898 253826 435454
rect 254382 434898 254414 435454
rect 253794 399454 254414 434898
rect 253794 398898 253826 399454
rect 254382 398898 254414 399454
rect 253794 363454 254414 398898
rect 253794 362898 253826 363454
rect 254382 362898 254414 363454
rect 253794 327454 254414 362898
rect 253794 326898 253826 327454
rect 254382 326898 254414 327454
rect 253794 291454 254414 326898
rect 253794 290898 253826 291454
rect 254382 290898 254414 291454
rect 253794 282628 254414 290898
rect 257514 705798 258134 711590
rect 257514 705242 257546 705798
rect 258102 705242 258134 705798
rect 257514 691174 258134 705242
rect 257514 690618 257546 691174
rect 258102 690618 258134 691174
rect 257514 655174 258134 690618
rect 257514 654618 257546 655174
rect 258102 654618 258134 655174
rect 257514 619174 258134 654618
rect 257514 618618 257546 619174
rect 258102 618618 258134 619174
rect 257514 583174 258134 618618
rect 257514 582618 257546 583174
rect 258102 582618 258134 583174
rect 257514 547174 258134 582618
rect 257514 546618 257546 547174
rect 258102 546618 258134 547174
rect 257514 511174 258134 546618
rect 257514 510618 257546 511174
rect 258102 510618 258134 511174
rect 257514 475174 258134 510618
rect 257514 474618 257546 475174
rect 258102 474618 258134 475174
rect 257514 439174 258134 474618
rect 257514 438618 257546 439174
rect 258102 438618 258134 439174
rect 257514 403174 258134 438618
rect 257514 402618 257546 403174
rect 258102 402618 258134 403174
rect 257514 367174 258134 402618
rect 257514 366618 257546 367174
rect 258102 366618 258134 367174
rect 257514 331174 258134 366618
rect 257514 330618 257546 331174
rect 258102 330618 258134 331174
rect 257514 295174 258134 330618
rect 257514 294618 257546 295174
rect 258102 294618 258134 295174
rect 243834 280938 243866 281494
rect 244422 280938 244454 281494
rect 243834 245494 244454 280938
rect 254288 274054 254608 274086
rect 254288 273818 254330 274054
rect 254566 273818 254608 274054
rect 254288 273734 254608 273818
rect 254288 273498 254330 273734
rect 254566 273498 254608 273734
rect 254288 273466 254608 273498
rect 246608 270334 246928 270366
rect 246608 270098 246650 270334
rect 246886 270098 246928 270334
rect 246608 270014 246928 270098
rect 246608 269778 246650 270014
rect 246886 269778 246928 270014
rect 246608 269746 246928 269778
rect 243834 244938 243866 245494
rect 244422 244938 244454 245494
rect 243834 209494 244454 244938
rect 257514 259174 258134 294618
rect 261234 706758 261854 711590
rect 261234 706202 261266 706758
rect 261822 706202 261854 706758
rect 261234 694894 261854 706202
rect 261234 694338 261266 694894
rect 261822 694338 261854 694894
rect 261234 658894 261854 694338
rect 261234 658338 261266 658894
rect 261822 658338 261854 658894
rect 261234 622894 261854 658338
rect 261234 622338 261266 622894
rect 261822 622338 261854 622894
rect 261234 586894 261854 622338
rect 261234 586338 261266 586894
rect 261822 586338 261854 586894
rect 261234 550894 261854 586338
rect 261234 550338 261266 550894
rect 261822 550338 261854 550894
rect 261234 514894 261854 550338
rect 261234 514338 261266 514894
rect 261822 514338 261854 514894
rect 261234 478894 261854 514338
rect 261234 478338 261266 478894
rect 261822 478338 261854 478894
rect 261234 442894 261854 478338
rect 261234 442338 261266 442894
rect 261822 442338 261854 442894
rect 261234 406894 261854 442338
rect 261234 406338 261266 406894
rect 261822 406338 261854 406894
rect 261234 370894 261854 406338
rect 261234 370338 261266 370894
rect 261822 370338 261854 370894
rect 261234 334894 261854 370338
rect 261234 334338 261266 334894
rect 261822 334338 261854 334894
rect 261234 298894 261854 334338
rect 261234 298338 261266 298894
rect 261822 298338 261854 298894
rect 261234 282628 261854 298338
rect 264954 707718 265574 711590
rect 264954 707162 264986 707718
rect 265542 707162 265574 707718
rect 264954 698614 265574 707162
rect 264954 698058 264986 698614
rect 265542 698058 265574 698614
rect 264954 662614 265574 698058
rect 264954 662058 264986 662614
rect 265542 662058 265574 662614
rect 264954 626614 265574 662058
rect 264954 626058 264986 626614
rect 265542 626058 265574 626614
rect 264954 590614 265574 626058
rect 264954 590058 264986 590614
rect 265542 590058 265574 590614
rect 264954 554614 265574 590058
rect 264954 554058 264986 554614
rect 265542 554058 265574 554614
rect 264954 518614 265574 554058
rect 264954 518058 264986 518614
rect 265542 518058 265574 518614
rect 264954 482614 265574 518058
rect 264954 482058 264986 482614
rect 265542 482058 265574 482614
rect 264954 446614 265574 482058
rect 264954 446058 264986 446614
rect 265542 446058 265574 446614
rect 264954 410614 265574 446058
rect 264954 410058 264986 410614
rect 265542 410058 265574 410614
rect 264954 374614 265574 410058
rect 264954 374058 264986 374614
rect 265542 374058 265574 374614
rect 264954 338614 265574 374058
rect 264954 338058 264986 338614
rect 265542 338058 265574 338614
rect 264954 302614 265574 338058
rect 264954 302058 264986 302614
rect 265542 302058 265574 302614
rect 257514 258618 257546 259174
rect 258102 258618 258134 259174
rect 254288 238054 254608 238086
rect 254288 237818 254330 238054
rect 254566 237818 254608 238054
rect 254288 237734 254608 237818
rect 254288 237498 254330 237734
rect 254566 237498 254608 237734
rect 254288 237466 254608 237498
rect 246608 234334 246928 234366
rect 246608 234098 246650 234334
rect 246886 234098 246928 234334
rect 246608 234014 246928 234098
rect 246608 233778 246650 234014
rect 246886 233778 246928 234014
rect 246608 233746 246928 233778
rect 243834 208938 243866 209494
rect 244422 208938 244454 209494
rect 243834 173494 244454 208938
rect 257514 223174 258134 258618
rect 264954 266614 265574 302058
rect 264954 266058 264986 266614
rect 265542 266058 265574 266614
rect 261968 255454 262288 255486
rect 261968 255218 262010 255454
rect 262246 255218 262288 255454
rect 261968 255134 262288 255218
rect 261968 254898 262010 255134
rect 262246 254898 262288 255134
rect 261968 254866 262288 254898
rect 257514 222618 257546 223174
rect 258102 222618 258134 223174
rect 254288 202054 254608 202086
rect 254288 201818 254330 202054
rect 254566 201818 254608 202054
rect 254288 201734 254608 201818
rect 254288 201498 254330 201734
rect 254566 201498 254608 201734
rect 254288 201466 254608 201498
rect 246608 198334 246928 198366
rect 246608 198098 246650 198334
rect 246886 198098 246928 198334
rect 246608 198014 246928 198098
rect 246608 197778 246650 198014
rect 246886 197778 246928 198014
rect 246608 197746 246928 197778
rect 243834 172938 243866 173494
rect 244422 172938 244454 173494
rect 243834 137494 244454 172938
rect 257514 187174 258134 222618
rect 264954 230614 265574 266058
rect 264954 230058 264986 230614
rect 265542 230058 265574 230614
rect 261968 219454 262288 219486
rect 261968 219218 262010 219454
rect 262246 219218 262288 219454
rect 261968 219134 262288 219218
rect 261968 218898 262010 219134
rect 262246 218898 262288 219134
rect 261968 218866 262288 218898
rect 257514 186618 257546 187174
rect 258102 186618 258134 187174
rect 254288 166054 254608 166086
rect 254288 165818 254330 166054
rect 254566 165818 254608 166054
rect 254288 165734 254608 165818
rect 254288 165498 254330 165734
rect 254566 165498 254608 165734
rect 254288 165466 254608 165498
rect 246608 162334 246928 162366
rect 246608 162098 246650 162334
rect 246886 162098 246928 162334
rect 246608 162014 246928 162098
rect 246608 161778 246650 162014
rect 246886 161778 246928 162014
rect 246608 161746 246928 161778
rect 243834 136938 243866 137494
rect 244422 136938 244454 137494
rect 243834 101494 244454 136938
rect 257514 151174 258134 186618
rect 264954 194614 265574 230058
rect 264954 194058 264986 194614
rect 265542 194058 265574 194614
rect 261968 183454 262288 183486
rect 261968 183218 262010 183454
rect 262246 183218 262288 183454
rect 261968 183134 262288 183218
rect 261968 182898 262010 183134
rect 262246 182898 262288 183134
rect 261968 182866 262288 182898
rect 257514 150618 257546 151174
rect 258102 150618 258134 151174
rect 254288 130054 254608 130086
rect 254288 129818 254330 130054
rect 254566 129818 254608 130054
rect 254288 129734 254608 129818
rect 254288 129498 254330 129734
rect 254566 129498 254608 129734
rect 254288 129466 254608 129498
rect 246608 126334 246928 126366
rect 246608 126098 246650 126334
rect 246886 126098 246928 126334
rect 246608 126014 246928 126098
rect 246608 125778 246650 126014
rect 246886 125778 246928 126014
rect 246608 125746 246928 125778
rect 243834 100938 243866 101494
rect 244422 100938 244454 101494
rect 243834 65494 244454 100938
rect 257514 115174 258134 150618
rect 264954 158614 265574 194058
rect 264954 158058 264986 158614
rect 265542 158058 265574 158614
rect 261968 147454 262288 147486
rect 261968 147218 262010 147454
rect 262246 147218 262288 147454
rect 261968 147134 262288 147218
rect 261968 146898 262010 147134
rect 262246 146898 262288 147134
rect 261968 146866 262288 146898
rect 257514 114618 257546 115174
rect 258102 114618 258134 115174
rect 254288 94054 254608 94086
rect 254288 93818 254330 94054
rect 254566 93818 254608 94054
rect 254288 93734 254608 93818
rect 254288 93498 254330 93734
rect 254566 93498 254608 93734
rect 254288 93466 254608 93498
rect 246608 90334 246928 90366
rect 246608 90098 246650 90334
rect 246886 90098 246928 90334
rect 246608 90014 246928 90098
rect 246608 89778 246650 90014
rect 246886 89778 246928 90014
rect 246608 89746 246928 89778
rect 243834 64938 243866 65494
rect 244422 64938 244454 65494
rect 243834 29494 244454 64938
rect 257514 79174 258134 114618
rect 264954 122614 265574 158058
rect 264954 122058 264986 122614
rect 265542 122058 265574 122614
rect 261968 111454 262288 111486
rect 261968 111218 262010 111454
rect 262246 111218 262288 111454
rect 261968 111134 262288 111218
rect 261968 110898 262010 111134
rect 262246 110898 262288 111134
rect 261968 110866 262288 110898
rect 257514 78618 257546 79174
rect 258102 78618 258134 79174
rect 254288 58054 254608 58086
rect 254288 57818 254330 58054
rect 254566 57818 254608 58054
rect 254288 57734 254608 57818
rect 254288 57498 254330 57734
rect 254566 57498 254608 57734
rect 254288 57466 254608 57498
rect 246608 54334 246928 54366
rect 246608 54098 246650 54334
rect 246886 54098 246928 54334
rect 246608 54014 246928 54098
rect 246608 53778 246650 54014
rect 246886 53778 246928 54014
rect 246608 53746 246928 53778
rect 243834 28938 243866 29494
rect 244422 28938 244454 29494
rect 243834 -7066 244454 28938
rect 257514 43174 258134 78618
rect 264954 86614 265574 122058
rect 264954 86058 264986 86614
rect 265542 86058 265574 86614
rect 261968 75454 262288 75486
rect 261968 75218 262010 75454
rect 262246 75218 262288 75454
rect 261968 75134 262288 75218
rect 261968 74898 262010 75134
rect 262246 74898 262288 75134
rect 261968 74866 262288 74898
rect 257514 42618 257546 43174
rect 258102 42618 258134 43174
rect 254288 22054 254608 22086
rect 254288 21818 254330 22054
rect 254566 21818 254608 22054
rect 254288 21734 254608 21818
rect 254288 21498 254330 21734
rect 254566 21498 254608 21734
rect 254288 21466 254608 21498
rect 246608 18334 246928 18366
rect 246608 18098 246650 18334
rect 246886 18098 246928 18334
rect 246608 18014 246928 18098
rect 246608 17778 246650 18014
rect 246886 17778 246928 18014
rect 246608 17746 246928 17778
rect 257514 7174 258134 42618
rect 264954 50614 265574 86058
rect 264954 50058 264986 50614
rect 265542 50058 265574 50614
rect 261968 39454 262288 39486
rect 261968 39218 262010 39454
rect 262246 39218 262288 39454
rect 261968 39134 262288 39218
rect 261968 38898 262010 39134
rect 262246 38898 262288 39134
rect 261968 38866 262288 38898
rect 257514 6618 257546 7174
rect 258102 6618 258134 7174
rect 243834 -7622 243866 -7066
rect 244422 -7622 244454 -7066
rect 243834 -7654 244454 -7622
rect 253794 -346 254414 2988
rect 253794 -902 253826 -346
rect 254382 -902 254414 -346
rect 253794 -7654 254414 -902
rect 257514 -1306 258134 6618
rect 264954 14614 265574 50058
rect 264954 14058 264986 14614
rect 265542 14058 265574 14614
rect 257514 -1862 257546 -1306
rect 258102 -1862 258134 -1306
rect 257514 -7654 258134 -1862
rect 261234 -2266 261854 2988
rect 261234 -2822 261266 -2266
rect 261822 -2822 261854 -2266
rect 261234 -7654 261854 -2822
rect 264954 -3226 265574 14058
rect 264954 -3782 264986 -3226
rect 265542 -3782 265574 -3226
rect 264954 -7654 265574 -3782
rect 268674 708678 269294 711590
rect 268674 708122 268706 708678
rect 269262 708122 269294 708678
rect 268674 666334 269294 708122
rect 268674 665778 268706 666334
rect 269262 665778 269294 666334
rect 268674 630334 269294 665778
rect 268674 629778 268706 630334
rect 269262 629778 269294 630334
rect 268674 594334 269294 629778
rect 268674 593778 268706 594334
rect 269262 593778 269294 594334
rect 268674 558334 269294 593778
rect 268674 557778 268706 558334
rect 269262 557778 269294 558334
rect 268674 522334 269294 557778
rect 268674 521778 268706 522334
rect 269262 521778 269294 522334
rect 268674 486334 269294 521778
rect 268674 485778 268706 486334
rect 269262 485778 269294 486334
rect 268674 450334 269294 485778
rect 268674 449778 268706 450334
rect 269262 449778 269294 450334
rect 268674 414334 269294 449778
rect 268674 413778 268706 414334
rect 269262 413778 269294 414334
rect 268674 378334 269294 413778
rect 268674 377778 268706 378334
rect 269262 377778 269294 378334
rect 268674 342334 269294 377778
rect 268674 341778 268706 342334
rect 269262 341778 269294 342334
rect 268674 306334 269294 341778
rect 268674 305778 268706 306334
rect 269262 305778 269294 306334
rect 268674 270334 269294 305778
rect 268674 269778 268706 270334
rect 269262 269778 269294 270334
rect 268674 234334 269294 269778
rect 272394 709638 273014 711590
rect 272394 709082 272426 709638
rect 272982 709082 273014 709638
rect 272394 670054 273014 709082
rect 272394 669498 272426 670054
rect 272982 669498 273014 670054
rect 272394 634054 273014 669498
rect 272394 633498 272426 634054
rect 272982 633498 273014 634054
rect 272394 598054 273014 633498
rect 272394 597498 272426 598054
rect 272982 597498 273014 598054
rect 272394 562054 273014 597498
rect 272394 561498 272426 562054
rect 272982 561498 273014 562054
rect 272394 526054 273014 561498
rect 272394 525498 272426 526054
rect 272982 525498 273014 526054
rect 272394 490054 273014 525498
rect 272394 489498 272426 490054
rect 272982 489498 273014 490054
rect 272394 454054 273014 489498
rect 272394 453498 272426 454054
rect 272982 453498 273014 454054
rect 272394 418054 273014 453498
rect 272394 417498 272426 418054
rect 272982 417498 273014 418054
rect 272394 382054 273014 417498
rect 272394 381498 272426 382054
rect 272982 381498 273014 382054
rect 272394 346054 273014 381498
rect 272394 345498 272426 346054
rect 272982 345498 273014 346054
rect 272394 310054 273014 345498
rect 272394 309498 272426 310054
rect 272982 309498 273014 310054
rect 272394 274054 273014 309498
rect 272394 273498 272426 274054
rect 272982 273498 273014 274054
rect 269648 259174 269968 259206
rect 269648 258938 269690 259174
rect 269926 258938 269968 259174
rect 269648 258854 269968 258938
rect 269648 258618 269690 258854
rect 269926 258618 269968 258854
rect 269648 258586 269968 258618
rect 268674 233778 268706 234334
rect 269262 233778 269294 234334
rect 268674 198334 269294 233778
rect 272394 238054 273014 273498
rect 272394 237498 272426 238054
rect 272982 237498 273014 238054
rect 269648 223174 269968 223206
rect 269648 222938 269690 223174
rect 269926 222938 269968 223174
rect 269648 222854 269968 222938
rect 269648 222618 269690 222854
rect 269926 222618 269968 222854
rect 269648 222586 269968 222618
rect 268674 197778 268706 198334
rect 269262 197778 269294 198334
rect 268674 162334 269294 197778
rect 272394 202054 273014 237498
rect 272394 201498 272426 202054
rect 272982 201498 273014 202054
rect 269648 187174 269968 187206
rect 269648 186938 269690 187174
rect 269926 186938 269968 187174
rect 269648 186854 269968 186938
rect 269648 186618 269690 186854
rect 269926 186618 269968 186854
rect 269648 186586 269968 186618
rect 268674 161778 268706 162334
rect 269262 161778 269294 162334
rect 268674 126334 269294 161778
rect 272394 166054 273014 201498
rect 272394 165498 272426 166054
rect 272982 165498 273014 166054
rect 269648 151174 269968 151206
rect 269648 150938 269690 151174
rect 269926 150938 269968 151174
rect 269648 150854 269968 150938
rect 269648 150618 269690 150854
rect 269926 150618 269968 150854
rect 269648 150586 269968 150618
rect 268674 125778 268706 126334
rect 269262 125778 269294 126334
rect 268674 90334 269294 125778
rect 272394 130054 273014 165498
rect 272394 129498 272426 130054
rect 272982 129498 273014 130054
rect 269648 115174 269968 115206
rect 269648 114938 269690 115174
rect 269926 114938 269968 115174
rect 269648 114854 269968 114938
rect 269648 114618 269690 114854
rect 269926 114618 269968 114854
rect 269648 114586 269968 114618
rect 268674 89778 268706 90334
rect 269262 89778 269294 90334
rect 268674 54334 269294 89778
rect 272394 94054 273014 129498
rect 272394 93498 272426 94054
rect 272982 93498 273014 94054
rect 269648 79174 269968 79206
rect 269648 78938 269690 79174
rect 269926 78938 269968 79174
rect 269648 78854 269968 78938
rect 269648 78618 269690 78854
rect 269926 78618 269968 78854
rect 269648 78586 269968 78618
rect 268674 53778 268706 54334
rect 269262 53778 269294 54334
rect 268674 18334 269294 53778
rect 272394 58054 273014 93498
rect 272394 57498 272426 58054
rect 272982 57498 273014 58054
rect 269648 43174 269968 43206
rect 269648 42938 269690 43174
rect 269926 42938 269968 43174
rect 269648 42854 269968 42938
rect 269648 42618 269690 42854
rect 269926 42618 269968 42854
rect 269648 42586 269968 42618
rect 268674 17778 268706 18334
rect 269262 17778 269294 18334
rect 268674 -4186 269294 17778
rect 272394 22054 273014 57498
rect 272394 21498 272426 22054
rect 272982 21498 273014 22054
rect 269648 7174 269968 7206
rect 269648 6938 269690 7174
rect 269926 6938 269968 7174
rect 269648 6854 269968 6938
rect 269648 6618 269690 6854
rect 269926 6618 269968 6854
rect 269648 6586 269968 6618
rect 268674 -4742 268706 -4186
rect 269262 -4742 269294 -4186
rect 268674 -7654 269294 -4742
rect 272394 -5146 273014 21498
rect 272394 -5702 272426 -5146
rect 272982 -5702 273014 -5146
rect 272394 -7654 273014 -5702
rect 276114 710598 276734 711590
rect 276114 710042 276146 710598
rect 276702 710042 276734 710598
rect 276114 673774 276734 710042
rect 276114 673218 276146 673774
rect 276702 673218 276734 673774
rect 276114 637774 276734 673218
rect 276114 637218 276146 637774
rect 276702 637218 276734 637774
rect 276114 601774 276734 637218
rect 276114 601218 276146 601774
rect 276702 601218 276734 601774
rect 276114 565774 276734 601218
rect 276114 565218 276146 565774
rect 276702 565218 276734 565774
rect 276114 529774 276734 565218
rect 276114 529218 276146 529774
rect 276702 529218 276734 529774
rect 276114 493774 276734 529218
rect 276114 493218 276146 493774
rect 276702 493218 276734 493774
rect 276114 457774 276734 493218
rect 276114 457218 276146 457774
rect 276702 457218 276734 457774
rect 276114 421774 276734 457218
rect 276114 421218 276146 421774
rect 276702 421218 276734 421774
rect 276114 385774 276734 421218
rect 276114 385218 276146 385774
rect 276702 385218 276734 385774
rect 276114 349774 276734 385218
rect 276114 349218 276146 349774
rect 276702 349218 276734 349774
rect 276114 313774 276734 349218
rect 276114 313218 276146 313774
rect 276702 313218 276734 313774
rect 276114 277774 276734 313218
rect 276114 277218 276146 277774
rect 276702 277218 276734 277774
rect 276114 241774 276734 277218
rect 279834 711558 280454 711590
rect 279834 711002 279866 711558
rect 280422 711002 280454 711558
rect 279834 677494 280454 711002
rect 279834 676938 279866 677494
rect 280422 676938 280454 677494
rect 279834 641494 280454 676938
rect 279834 640938 279866 641494
rect 280422 640938 280454 641494
rect 279834 605494 280454 640938
rect 279834 604938 279866 605494
rect 280422 604938 280454 605494
rect 279834 569494 280454 604938
rect 279834 568938 279866 569494
rect 280422 568938 280454 569494
rect 279834 533494 280454 568938
rect 279834 532938 279866 533494
rect 280422 532938 280454 533494
rect 279834 497494 280454 532938
rect 279834 496938 279866 497494
rect 280422 496938 280454 497494
rect 279834 461494 280454 496938
rect 279834 460938 279866 461494
rect 280422 460938 280454 461494
rect 279834 425494 280454 460938
rect 279834 424938 279866 425494
rect 280422 424938 280454 425494
rect 279834 389494 280454 424938
rect 279834 388938 279866 389494
rect 280422 388938 280454 389494
rect 279834 353494 280454 388938
rect 279834 352938 279866 353494
rect 280422 352938 280454 353494
rect 279834 317494 280454 352938
rect 279834 316938 279866 317494
rect 280422 316938 280454 317494
rect 279834 281494 280454 316938
rect 279834 280938 279866 281494
rect 280422 280938 280454 281494
rect 277328 270334 277648 270366
rect 277328 270098 277370 270334
rect 277606 270098 277648 270334
rect 277328 270014 277648 270098
rect 277328 269778 277370 270014
rect 277606 269778 277648 270014
rect 277328 269746 277648 269778
rect 276114 241218 276146 241774
rect 276702 241218 276734 241774
rect 276114 205774 276734 241218
rect 279834 245494 280454 280938
rect 289794 704838 290414 711590
rect 289794 704282 289826 704838
rect 290382 704282 290414 704838
rect 289794 687454 290414 704282
rect 289794 686898 289826 687454
rect 290382 686898 290414 687454
rect 289794 651454 290414 686898
rect 289794 650898 289826 651454
rect 290382 650898 290414 651454
rect 289794 615454 290414 650898
rect 289794 614898 289826 615454
rect 290382 614898 290414 615454
rect 289794 579454 290414 614898
rect 289794 578898 289826 579454
rect 290382 578898 290414 579454
rect 289794 543454 290414 578898
rect 289794 542898 289826 543454
rect 290382 542898 290414 543454
rect 289794 507454 290414 542898
rect 289794 506898 289826 507454
rect 290382 506898 290414 507454
rect 289794 471454 290414 506898
rect 289794 470898 289826 471454
rect 290382 470898 290414 471454
rect 289794 435454 290414 470898
rect 289794 434898 289826 435454
rect 290382 434898 290414 435454
rect 289794 399454 290414 434898
rect 289794 398898 289826 399454
rect 290382 398898 290414 399454
rect 289794 363454 290414 398898
rect 289794 362898 289826 363454
rect 290382 362898 290414 363454
rect 289794 327454 290414 362898
rect 289794 326898 289826 327454
rect 290382 326898 290414 327454
rect 289794 291454 290414 326898
rect 289794 290898 289826 291454
rect 290382 290898 290414 291454
rect 285008 274054 285328 274086
rect 285008 273818 285050 274054
rect 285286 273818 285328 274054
rect 285008 273734 285328 273818
rect 285008 273498 285050 273734
rect 285286 273498 285328 273734
rect 285008 273466 285328 273498
rect 279834 244938 279866 245494
rect 280422 244938 280454 245494
rect 277328 234334 277648 234366
rect 277328 234098 277370 234334
rect 277606 234098 277648 234334
rect 277328 234014 277648 234098
rect 277328 233778 277370 234014
rect 277606 233778 277648 234014
rect 277328 233746 277648 233778
rect 276114 205218 276146 205774
rect 276702 205218 276734 205774
rect 276114 169774 276734 205218
rect 279834 209494 280454 244938
rect 289794 255454 290414 290898
rect 289794 254898 289826 255454
rect 290382 254898 290414 255454
rect 285008 238054 285328 238086
rect 285008 237818 285050 238054
rect 285286 237818 285328 238054
rect 285008 237734 285328 237818
rect 285008 237498 285050 237734
rect 285286 237498 285328 237734
rect 285008 237466 285328 237498
rect 279834 208938 279866 209494
rect 280422 208938 280454 209494
rect 277328 198334 277648 198366
rect 277328 198098 277370 198334
rect 277606 198098 277648 198334
rect 277328 198014 277648 198098
rect 277328 197778 277370 198014
rect 277606 197778 277648 198014
rect 277328 197746 277648 197778
rect 276114 169218 276146 169774
rect 276702 169218 276734 169774
rect 276114 133774 276734 169218
rect 279834 173494 280454 208938
rect 289794 219454 290414 254898
rect 289794 218898 289826 219454
rect 290382 218898 290414 219454
rect 285008 202054 285328 202086
rect 285008 201818 285050 202054
rect 285286 201818 285328 202054
rect 285008 201734 285328 201818
rect 285008 201498 285050 201734
rect 285286 201498 285328 201734
rect 285008 201466 285328 201498
rect 279834 172938 279866 173494
rect 280422 172938 280454 173494
rect 277328 162334 277648 162366
rect 277328 162098 277370 162334
rect 277606 162098 277648 162334
rect 277328 162014 277648 162098
rect 277328 161778 277370 162014
rect 277606 161778 277648 162014
rect 277328 161746 277648 161778
rect 276114 133218 276146 133774
rect 276702 133218 276734 133774
rect 276114 97774 276734 133218
rect 279834 137494 280454 172938
rect 289794 183454 290414 218898
rect 289794 182898 289826 183454
rect 290382 182898 290414 183454
rect 285008 166054 285328 166086
rect 285008 165818 285050 166054
rect 285286 165818 285328 166054
rect 285008 165734 285328 165818
rect 285008 165498 285050 165734
rect 285286 165498 285328 165734
rect 285008 165466 285328 165498
rect 279834 136938 279866 137494
rect 280422 136938 280454 137494
rect 277328 126334 277648 126366
rect 277328 126098 277370 126334
rect 277606 126098 277648 126334
rect 277328 126014 277648 126098
rect 277328 125778 277370 126014
rect 277606 125778 277648 126014
rect 277328 125746 277648 125778
rect 276114 97218 276146 97774
rect 276702 97218 276734 97774
rect 276114 61774 276734 97218
rect 279834 101494 280454 136938
rect 289794 147454 290414 182898
rect 289794 146898 289826 147454
rect 290382 146898 290414 147454
rect 285008 130054 285328 130086
rect 285008 129818 285050 130054
rect 285286 129818 285328 130054
rect 285008 129734 285328 129818
rect 285008 129498 285050 129734
rect 285286 129498 285328 129734
rect 285008 129466 285328 129498
rect 279834 100938 279866 101494
rect 280422 100938 280454 101494
rect 277328 90334 277648 90366
rect 277328 90098 277370 90334
rect 277606 90098 277648 90334
rect 277328 90014 277648 90098
rect 277328 89778 277370 90014
rect 277606 89778 277648 90014
rect 277328 89746 277648 89778
rect 276114 61218 276146 61774
rect 276702 61218 276734 61774
rect 276114 25774 276734 61218
rect 279834 65494 280454 100938
rect 289794 111454 290414 146898
rect 289794 110898 289826 111454
rect 290382 110898 290414 111454
rect 285008 94054 285328 94086
rect 285008 93818 285050 94054
rect 285286 93818 285328 94054
rect 285008 93734 285328 93818
rect 285008 93498 285050 93734
rect 285286 93498 285328 93734
rect 285008 93466 285328 93498
rect 279834 64938 279866 65494
rect 280422 64938 280454 65494
rect 277328 54334 277648 54366
rect 277328 54098 277370 54334
rect 277606 54098 277648 54334
rect 277328 54014 277648 54098
rect 277328 53778 277370 54014
rect 277606 53778 277648 54014
rect 277328 53746 277648 53778
rect 276114 25218 276146 25774
rect 276702 25218 276734 25774
rect 276114 -6106 276734 25218
rect 279834 29494 280454 64938
rect 289794 75454 290414 110898
rect 289794 74898 289826 75454
rect 290382 74898 290414 75454
rect 285008 58054 285328 58086
rect 285008 57818 285050 58054
rect 285286 57818 285328 58054
rect 285008 57734 285328 57818
rect 285008 57498 285050 57734
rect 285286 57498 285328 57734
rect 285008 57466 285328 57498
rect 279834 28938 279866 29494
rect 280422 28938 280454 29494
rect 277328 18334 277648 18366
rect 277328 18098 277370 18334
rect 277606 18098 277648 18334
rect 277328 18014 277648 18098
rect 277328 17778 277370 18014
rect 277606 17778 277648 18014
rect 277328 17746 277648 17778
rect 276114 -6662 276146 -6106
rect 276702 -6662 276734 -6106
rect 276114 -7654 276734 -6662
rect 279834 -7066 280454 28938
rect 289794 39454 290414 74898
rect 289794 38898 289826 39454
rect 290382 38898 290414 39454
rect 285008 22054 285328 22086
rect 285008 21818 285050 22054
rect 285286 21818 285328 22054
rect 285008 21734 285328 21818
rect 285008 21498 285050 21734
rect 285286 21498 285328 21734
rect 285008 21466 285328 21498
rect 279834 -7622 279866 -7066
rect 280422 -7622 280454 -7066
rect 279834 -7654 280454 -7622
rect 289794 3454 290414 38898
rect 289794 2898 289826 3454
rect 290382 2898 290414 3454
rect 289794 -346 290414 2898
rect 289794 -902 289826 -346
rect 290382 -902 290414 -346
rect 289794 -7654 290414 -902
rect 293514 705798 294134 711590
rect 293514 705242 293546 705798
rect 294102 705242 294134 705798
rect 293514 691174 294134 705242
rect 293514 690618 293546 691174
rect 294102 690618 294134 691174
rect 293514 655174 294134 690618
rect 293514 654618 293546 655174
rect 294102 654618 294134 655174
rect 293514 619174 294134 654618
rect 293514 618618 293546 619174
rect 294102 618618 294134 619174
rect 293514 583174 294134 618618
rect 293514 582618 293546 583174
rect 294102 582618 294134 583174
rect 293514 547174 294134 582618
rect 293514 546618 293546 547174
rect 294102 546618 294134 547174
rect 293514 511174 294134 546618
rect 293514 510618 293546 511174
rect 294102 510618 294134 511174
rect 293514 475174 294134 510618
rect 293514 474618 293546 475174
rect 294102 474618 294134 475174
rect 293514 439174 294134 474618
rect 293514 438618 293546 439174
rect 294102 438618 294134 439174
rect 293514 403174 294134 438618
rect 293514 402618 293546 403174
rect 294102 402618 294134 403174
rect 293514 367174 294134 402618
rect 293514 366618 293546 367174
rect 294102 366618 294134 367174
rect 293514 331174 294134 366618
rect 293514 330618 293546 331174
rect 294102 330618 294134 331174
rect 293514 295174 294134 330618
rect 293514 294618 293546 295174
rect 294102 294618 294134 295174
rect 293514 259174 294134 294618
rect 293514 258618 293546 259174
rect 294102 258618 294134 259174
rect 293514 223174 294134 258618
rect 293514 222618 293546 223174
rect 294102 222618 294134 223174
rect 293514 187174 294134 222618
rect 293514 186618 293546 187174
rect 294102 186618 294134 187174
rect 293514 151174 294134 186618
rect 293514 150618 293546 151174
rect 294102 150618 294134 151174
rect 293514 115174 294134 150618
rect 293514 114618 293546 115174
rect 294102 114618 294134 115174
rect 293514 79174 294134 114618
rect 293514 78618 293546 79174
rect 294102 78618 294134 79174
rect 293514 43174 294134 78618
rect 293514 42618 293546 43174
rect 294102 42618 294134 43174
rect 293514 7174 294134 42618
rect 293514 6618 293546 7174
rect 294102 6618 294134 7174
rect 293514 -1306 294134 6618
rect 293514 -1862 293546 -1306
rect 294102 -1862 294134 -1306
rect 293514 -7654 294134 -1862
rect 297234 706758 297854 711590
rect 297234 706202 297266 706758
rect 297822 706202 297854 706758
rect 297234 694894 297854 706202
rect 297234 694338 297266 694894
rect 297822 694338 297854 694894
rect 297234 658894 297854 694338
rect 297234 658338 297266 658894
rect 297822 658338 297854 658894
rect 297234 622894 297854 658338
rect 297234 622338 297266 622894
rect 297822 622338 297854 622894
rect 297234 586894 297854 622338
rect 297234 586338 297266 586894
rect 297822 586338 297854 586894
rect 297234 550894 297854 586338
rect 297234 550338 297266 550894
rect 297822 550338 297854 550894
rect 297234 514894 297854 550338
rect 297234 514338 297266 514894
rect 297822 514338 297854 514894
rect 297234 478894 297854 514338
rect 297234 478338 297266 478894
rect 297822 478338 297854 478894
rect 297234 442894 297854 478338
rect 297234 442338 297266 442894
rect 297822 442338 297854 442894
rect 297234 406894 297854 442338
rect 297234 406338 297266 406894
rect 297822 406338 297854 406894
rect 297234 370894 297854 406338
rect 297234 370338 297266 370894
rect 297822 370338 297854 370894
rect 297234 334894 297854 370338
rect 297234 334338 297266 334894
rect 297822 334338 297854 334894
rect 297234 298894 297854 334338
rect 297234 298338 297266 298894
rect 297822 298338 297854 298894
rect 297234 262894 297854 298338
rect 297234 262338 297266 262894
rect 297822 262338 297854 262894
rect 297234 226894 297854 262338
rect 297234 226338 297266 226894
rect 297822 226338 297854 226894
rect 297234 190894 297854 226338
rect 297234 190338 297266 190894
rect 297822 190338 297854 190894
rect 297234 154894 297854 190338
rect 297234 154338 297266 154894
rect 297822 154338 297854 154894
rect 297234 118894 297854 154338
rect 297234 118338 297266 118894
rect 297822 118338 297854 118894
rect 297234 82894 297854 118338
rect 297234 82338 297266 82894
rect 297822 82338 297854 82894
rect 297234 46894 297854 82338
rect 297234 46338 297266 46894
rect 297822 46338 297854 46894
rect 297234 10894 297854 46338
rect 297234 10338 297266 10894
rect 297822 10338 297854 10894
rect 297234 -2266 297854 10338
rect 297234 -2822 297266 -2266
rect 297822 -2822 297854 -2266
rect 297234 -7654 297854 -2822
rect 300954 707718 301574 711590
rect 300954 707162 300986 707718
rect 301542 707162 301574 707718
rect 300954 698614 301574 707162
rect 300954 698058 300986 698614
rect 301542 698058 301574 698614
rect 300954 662614 301574 698058
rect 300954 662058 300986 662614
rect 301542 662058 301574 662614
rect 300954 626614 301574 662058
rect 300954 626058 300986 626614
rect 301542 626058 301574 626614
rect 300954 590614 301574 626058
rect 300954 590058 300986 590614
rect 301542 590058 301574 590614
rect 300954 554614 301574 590058
rect 300954 554058 300986 554614
rect 301542 554058 301574 554614
rect 300954 518614 301574 554058
rect 300954 518058 300986 518614
rect 301542 518058 301574 518614
rect 300954 482614 301574 518058
rect 300954 482058 300986 482614
rect 301542 482058 301574 482614
rect 300954 446614 301574 482058
rect 300954 446058 300986 446614
rect 301542 446058 301574 446614
rect 300954 410614 301574 446058
rect 300954 410058 300986 410614
rect 301542 410058 301574 410614
rect 300954 374614 301574 410058
rect 300954 374058 300986 374614
rect 301542 374058 301574 374614
rect 300954 338614 301574 374058
rect 300954 338058 300986 338614
rect 301542 338058 301574 338614
rect 300954 302614 301574 338058
rect 300954 302058 300986 302614
rect 301542 302058 301574 302614
rect 300954 266614 301574 302058
rect 300954 266058 300986 266614
rect 301542 266058 301574 266614
rect 300954 230614 301574 266058
rect 300954 230058 300986 230614
rect 301542 230058 301574 230614
rect 300954 194614 301574 230058
rect 300954 194058 300986 194614
rect 301542 194058 301574 194614
rect 300954 158614 301574 194058
rect 300954 158058 300986 158614
rect 301542 158058 301574 158614
rect 300954 122614 301574 158058
rect 300954 122058 300986 122614
rect 301542 122058 301574 122614
rect 300954 86614 301574 122058
rect 300954 86058 300986 86614
rect 301542 86058 301574 86614
rect 300954 50614 301574 86058
rect 300954 50058 300986 50614
rect 301542 50058 301574 50614
rect 300954 14614 301574 50058
rect 300954 14058 300986 14614
rect 301542 14058 301574 14614
rect 300954 -3226 301574 14058
rect 300954 -3782 300986 -3226
rect 301542 -3782 301574 -3226
rect 300954 -7654 301574 -3782
rect 304674 708678 305294 711590
rect 304674 708122 304706 708678
rect 305262 708122 305294 708678
rect 304674 666334 305294 708122
rect 304674 665778 304706 666334
rect 305262 665778 305294 666334
rect 304674 630334 305294 665778
rect 304674 629778 304706 630334
rect 305262 629778 305294 630334
rect 304674 594334 305294 629778
rect 304674 593778 304706 594334
rect 305262 593778 305294 594334
rect 304674 558334 305294 593778
rect 304674 557778 304706 558334
rect 305262 557778 305294 558334
rect 304674 522334 305294 557778
rect 304674 521778 304706 522334
rect 305262 521778 305294 522334
rect 304674 486334 305294 521778
rect 304674 485778 304706 486334
rect 305262 485778 305294 486334
rect 304674 450334 305294 485778
rect 304674 449778 304706 450334
rect 305262 449778 305294 450334
rect 304674 414334 305294 449778
rect 304674 413778 304706 414334
rect 305262 413778 305294 414334
rect 304674 378334 305294 413778
rect 304674 377778 304706 378334
rect 305262 377778 305294 378334
rect 304674 342334 305294 377778
rect 304674 341778 304706 342334
rect 305262 341778 305294 342334
rect 304674 306334 305294 341778
rect 304674 305778 304706 306334
rect 305262 305778 305294 306334
rect 304674 270334 305294 305778
rect 304674 269778 304706 270334
rect 305262 269778 305294 270334
rect 304674 234334 305294 269778
rect 304674 233778 304706 234334
rect 305262 233778 305294 234334
rect 304674 198334 305294 233778
rect 304674 197778 304706 198334
rect 305262 197778 305294 198334
rect 304674 162334 305294 197778
rect 304674 161778 304706 162334
rect 305262 161778 305294 162334
rect 304674 126334 305294 161778
rect 304674 125778 304706 126334
rect 305262 125778 305294 126334
rect 304674 90334 305294 125778
rect 304674 89778 304706 90334
rect 305262 89778 305294 90334
rect 304674 54334 305294 89778
rect 304674 53778 304706 54334
rect 305262 53778 305294 54334
rect 304674 18334 305294 53778
rect 304674 17778 304706 18334
rect 305262 17778 305294 18334
rect 304674 -4186 305294 17778
rect 304674 -4742 304706 -4186
rect 305262 -4742 305294 -4186
rect 304674 -7654 305294 -4742
rect 308394 709638 309014 711590
rect 308394 709082 308426 709638
rect 308982 709082 309014 709638
rect 308394 670054 309014 709082
rect 308394 669498 308426 670054
rect 308982 669498 309014 670054
rect 308394 634054 309014 669498
rect 308394 633498 308426 634054
rect 308982 633498 309014 634054
rect 308394 598054 309014 633498
rect 308394 597498 308426 598054
rect 308982 597498 309014 598054
rect 308394 562054 309014 597498
rect 308394 561498 308426 562054
rect 308982 561498 309014 562054
rect 308394 526054 309014 561498
rect 308394 525498 308426 526054
rect 308982 525498 309014 526054
rect 308394 490054 309014 525498
rect 308394 489498 308426 490054
rect 308982 489498 309014 490054
rect 308394 454054 309014 489498
rect 308394 453498 308426 454054
rect 308982 453498 309014 454054
rect 308394 418054 309014 453498
rect 308394 417498 308426 418054
rect 308982 417498 309014 418054
rect 308394 382054 309014 417498
rect 308394 381498 308426 382054
rect 308982 381498 309014 382054
rect 308394 346054 309014 381498
rect 308394 345498 308426 346054
rect 308982 345498 309014 346054
rect 308394 310054 309014 345498
rect 308394 309498 308426 310054
rect 308982 309498 309014 310054
rect 308394 274054 309014 309498
rect 308394 273498 308426 274054
rect 308982 273498 309014 274054
rect 308394 238054 309014 273498
rect 308394 237498 308426 238054
rect 308982 237498 309014 238054
rect 308394 202054 309014 237498
rect 308394 201498 308426 202054
rect 308982 201498 309014 202054
rect 308394 166054 309014 201498
rect 308394 165498 308426 166054
rect 308982 165498 309014 166054
rect 308394 130054 309014 165498
rect 308394 129498 308426 130054
rect 308982 129498 309014 130054
rect 308394 94054 309014 129498
rect 308394 93498 308426 94054
rect 308982 93498 309014 94054
rect 308394 58054 309014 93498
rect 308394 57498 308426 58054
rect 308982 57498 309014 58054
rect 308394 22054 309014 57498
rect 308394 21498 308426 22054
rect 308982 21498 309014 22054
rect 308394 -5146 309014 21498
rect 308394 -5702 308426 -5146
rect 308982 -5702 309014 -5146
rect 308394 -7654 309014 -5702
rect 312114 710598 312734 711590
rect 312114 710042 312146 710598
rect 312702 710042 312734 710598
rect 312114 673774 312734 710042
rect 312114 673218 312146 673774
rect 312702 673218 312734 673774
rect 312114 637774 312734 673218
rect 312114 637218 312146 637774
rect 312702 637218 312734 637774
rect 312114 601774 312734 637218
rect 312114 601218 312146 601774
rect 312702 601218 312734 601774
rect 312114 565774 312734 601218
rect 312114 565218 312146 565774
rect 312702 565218 312734 565774
rect 312114 529774 312734 565218
rect 312114 529218 312146 529774
rect 312702 529218 312734 529774
rect 312114 493774 312734 529218
rect 312114 493218 312146 493774
rect 312702 493218 312734 493774
rect 312114 457774 312734 493218
rect 312114 457218 312146 457774
rect 312702 457218 312734 457774
rect 312114 421774 312734 457218
rect 312114 421218 312146 421774
rect 312702 421218 312734 421774
rect 312114 385774 312734 421218
rect 312114 385218 312146 385774
rect 312702 385218 312734 385774
rect 312114 349774 312734 385218
rect 312114 349218 312146 349774
rect 312702 349218 312734 349774
rect 312114 313774 312734 349218
rect 312114 313218 312146 313774
rect 312702 313218 312734 313774
rect 312114 277774 312734 313218
rect 312114 277218 312146 277774
rect 312702 277218 312734 277774
rect 312114 241774 312734 277218
rect 312114 241218 312146 241774
rect 312702 241218 312734 241774
rect 312114 205774 312734 241218
rect 312114 205218 312146 205774
rect 312702 205218 312734 205774
rect 312114 169774 312734 205218
rect 312114 169218 312146 169774
rect 312702 169218 312734 169774
rect 312114 133774 312734 169218
rect 312114 133218 312146 133774
rect 312702 133218 312734 133774
rect 312114 97774 312734 133218
rect 312114 97218 312146 97774
rect 312702 97218 312734 97774
rect 312114 61774 312734 97218
rect 312114 61218 312146 61774
rect 312702 61218 312734 61774
rect 312114 25774 312734 61218
rect 312114 25218 312146 25774
rect 312702 25218 312734 25774
rect 312114 -6106 312734 25218
rect 312114 -6662 312146 -6106
rect 312702 -6662 312734 -6106
rect 312114 -7654 312734 -6662
rect 315834 711558 316454 711590
rect 315834 711002 315866 711558
rect 316422 711002 316454 711558
rect 315834 677494 316454 711002
rect 315834 676938 315866 677494
rect 316422 676938 316454 677494
rect 315834 641494 316454 676938
rect 315834 640938 315866 641494
rect 316422 640938 316454 641494
rect 315834 605494 316454 640938
rect 315834 604938 315866 605494
rect 316422 604938 316454 605494
rect 315834 569494 316454 604938
rect 315834 568938 315866 569494
rect 316422 568938 316454 569494
rect 315834 533494 316454 568938
rect 315834 532938 315866 533494
rect 316422 532938 316454 533494
rect 315834 497494 316454 532938
rect 315834 496938 315866 497494
rect 316422 496938 316454 497494
rect 315834 461494 316454 496938
rect 315834 460938 315866 461494
rect 316422 460938 316454 461494
rect 315834 425494 316454 460938
rect 315834 424938 315866 425494
rect 316422 424938 316454 425494
rect 315834 389494 316454 424938
rect 315834 388938 315866 389494
rect 316422 388938 316454 389494
rect 315834 353494 316454 388938
rect 315834 352938 315866 353494
rect 316422 352938 316454 353494
rect 315834 317494 316454 352938
rect 315834 316938 315866 317494
rect 316422 316938 316454 317494
rect 315834 281494 316454 316938
rect 315834 280938 315866 281494
rect 316422 280938 316454 281494
rect 315834 245494 316454 280938
rect 315834 244938 315866 245494
rect 316422 244938 316454 245494
rect 315834 209494 316454 244938
rect 315834 208938 315866 209494
rect 316422 208938 316454 209494
rect 315834 173494 316454 208938
rect 315834 172938 315866 173494
rect 316422 172938 316454 173494
rect 315834 137494 316454 172938
rect 315834 136938 315866 137494
rect 316422 136938 316454 137494
rect 315834 101494 316454 136938
rect 315834 100938 315866 101494
rect 316422 100938 316454 101494
rect 315834 65494 316454 100938
rect 315834 64938 315866 65494
rect 316422 64938 316454 65494
rect 315834 29494 316454 64938
rect 315834 28938 315866 29494
rect 316422 28938 316454 29494
rect 315834 -7066 316454 28938
rect 315834 -7622 315866 -7066
rect 316422 -7622 316454 -7066
rect 315834 -7654 316454 -7622
rect 325794 704838 326414 711590
rect 325794 704282 325826 704838
rect 326382 704282 326414 704838
rect 325794 687454 326414 704282
rect 325794 686898 325826 687454
rect 326382 686898 326414 687454
rect 325794 651454 326414 686898
rect 325794 650898 325826 651454
rect 326382 650898 326414 651454
rect 325794 615454 326414 650898
rect 325794 614898 325826 615454
rect 326382 614898 326414 615454
rect 325794 579454 326414 614898
rect 325794 578898 325826 579454
rect 326382 578898 326414 579454
rect 325794 543454 326414 578898
rect 325794 542898 325826 543454
rect 326382 542898 326414 543454
rect 325794 507454 326414 542898
rect 325794 506898 325826 507454
rect 326382 506898 326414 507454
rect 325794 471454 326414 506898
rect 325794 470898 325826 471454
rect 326382 470898 326414 471454
rect 325794 435454 326414 470898
rect 325794 434898 325826 435454
rect 326382 434898 326414 435454
rect 325794 399454 326414 434898
rect 325794 398898 325826 399454
rect 326382 398898 326414 399454
rect 325794 363454 326414 398898
rect 325794 362898 325826 363454
rect 326382 362898 326414 363454
rect 325794 327454 326414 362898
rect 325794 326898 325826 327454
rect 326382 326898 326414 327454
rect 325794 291454 326414 326898
rect 325794 290898 325826 291454
rect 326382 290898 326414 291454
rect 325794 255454 326414 290898
rect 325794 254898 325826 255454
rect 326382 254898 326414 255454
rect 325794 219454 326414 254898
rect 325794 218898 325826 219454
rect 326382 218898 326414 219454
rect 325794 183454 326414 218898
rect 325794 182898 325826 183454
rect 326382 182898 326414 183454
rect 325794 147454 326414 182898
rect 325794 146898 325826 147454
rect 326382 146898 326414 147454
rect 325794 111454 326414 146898
rect 325794 110898 325826 111454
rect 326382 110898 326414 111454
rect 325794 75454 326414 110898
rect 325794 74898 325826 75454
rect 326382 74898 326414 75454
rect 325794 39454 326414 74898
rect 325794 38898 325826 39454
rect 326382 38898 326414 39454
rect 325794 3454 326414 38898
rect 325794 2898 325826 3454
rect 326382 2898 326414 3454
rect 325794 -346 326414 2898
rect 325794 -902 325826 -346
rect 326382 -902 326414 -346
rect 325794 -7654 326414 -902
rect 329514 705798 330134 711590
rect 329514 705242 329546 705798
rect 330102 705242 330134 705798
rect 329514 691174 330134 705242
rect 329514 690618 329546 691174
rect 330102 690618 330134 691174
rect 329514 655174 330134 690618
rect 329514 654618 329546 655174
rect 330102 654618 330134 655174
rect 329514 619174 330134 654618
rect 329514 618618 329546 619174
rect 330102 618618 330134 619174
rect 329514 583174 330134 618618
rect 329514 582618 329546 583174
rect 330102 582618 330134 583174
rect 329514 547174 330134 582618
rect 329514 546618 329546 547174
rect 330102 546618 330134 547174
rect 329514 511174 330134 546618
rect 329514 510618 329546 511174
rect 330102 510618 330134 511174
rect 329514 475174 330134 510618
rect 329514 474618 329546 475174
rect 330102 474618 330134 475174
rect 329514 439174 330134 474618
rect 329514 438618 329546 439174
rect 330102 438618 330134 439174
rect 329514 403174 330134 438618
rect 329514 402618 329546 403174
rect 330102 402618 330134 403174
rect 329514 367174 330134 402618
rect 329514 366618 329546 367174
rect 330102 366618 330134 367174
rect 329514 331174 330134 366618
rect 329514 330618 329546 331174
rect 330102 330618 330134 331174
rect 329514 295174 330134 330618
rect 329514 294618 329546 295174
rect 330102 294618 330134 295174
rect 329514 259174 330134 294618
rect 329514 258618 329546 259174
rect 330102 258618 330134 259174
rect 329514 223174 330134 258618
rect 329514 222618 329546 223174
rect 330102 222618 330134 223174
rect 329514 187174 330134 222618
rect 329514 186618 329546 187174
rect 330102 186618 330134 187174
rect 329514 151174 330134 186618
rect 329514 150618 329546 151174
rect 330102 150618 330134 151174
rect 329514 115174 330134 150618
rect 329514 114618 329546 115174
rect 330102 114618 330134 115174
rect 329514 79174 330134 114618
rect 329514 78618 329546 79174
rect 330102 78618 330134 79174
rect 329514 43174 330134 78618
rect 329514 42618 329546 43174
rect 330102 42618 330134 43174
rect 329514 7174 330134 42618
rect 329514 6618 329546 7174
rect 330102 6618 330134 7174
rect 329514 -1306 330134 6618
rect 329514 -1862 329546 -1306
rect 330102 -1862 330134 -1306
rect 329514 -7654 330134 -1862
rect 333234 706758 333854 711590
rect 333234 706202 333266 706758
rect 333822 706202 333854 706758
rect 333234 694894 333854 706202
rect 333234 694338 333266 694894
rect 333822 694338 333854 694894
rect 333234 658894 333854 694338
rect 333234 658338 333266 658894
rect 333822 658338 333854 658894
rect 333234 622894 333854 658338
rect 333234 622338 333266 622894
rect 333822 622338 333854 622894
rect 333234 586894 333854 622338
rect 333234 586338 333266 586894
rect 333822 586338 333854 586894
rect 333234 550894 333854 586338
rect 333234 550338 333266 550894
rect 333822 550338 333854 550894
rect 333234 514894 333854 550338
rect 333234 514338 333266 514894
rect 333822 514338 333854 514894
rect 333234 478894 333854 514338
rect 333234 478338 333266 478894
rect 333822 478338 333854 478894
rect 333234 442894 333854 478338
rect 333234 442338 333266 442894
rect 333822 442338 333854 442894
rect 333234 406894 333854 442338
rect 333234 406338 333266 406894
rect 333822 406338 333854 406894
rect 333234 370894 333854 406338
rect 333234 370338 333266 370894
rect 333822 370338 333854 370894
rect 333234 334894 333854 370338
rect 333234 334338 333266 334894
rect 333822 334338 333854 334894
rect 333234 298894 333854 334338
rect 333234 298338 333266 298894
rect 333822 298338 333854 298894
rect 333234 262894 333854 298338
rect 333234 262338 333266 262894
rect 333822 262338 333854 262894
rect 333234 226894 333854 262338
rect 333234 226338 333266 226894
rect 333822 226338 333854 226894
rect 333234 190894 333854 226338
rect 333234 190338 333266 190894
rect 333822 190338 333854 190894
rect 333234 154894 333854 190338
rect 333234 154338 333266 154894
rect 333822 154338 333854 154894
rect 333234 118894 333854 154338
rect 333234 118338 333266 118894
rect 333822 118338 333854 118894
rect 333234 82894 333854 118338
rect 333234 82338 333266 82894
rect 333822 82338 333854 82894
rect 333234 46894 333854 82338
rect 333234 46338 333266 46894
rect 333822 46338 333854 46894
rect 333234 10894 333854 46338
rect 333234 10338 333266 10894
rect 333822 10338 333854 10894
rect 333234 -2266 333854 10338
rect 333234 -2822 333266 -2266
rect 333822 -2822 333854 -2266
rect 333234 -7654 333854 -2822
rect 336954 707718 337574 711590
rect 336954 707162 336986 707718
rect 337542 707162 337574 707718
rect 336954 698614 337574 707162
rect 336954 698058 336986 698614
rect 337542 698058 337574 698614
rect 336954 662614 337574 698058
rect 336954 662058 336986 662614
rect 337542 662058 337574 662614
rect 336954 626614 337574 662058
rect 336954 626058 336986 626614
rect 337542 626058 337574 626614
rect 336954 590614 337574 626058
rect 336954 590058 336986 590614
rect 337542 590058 337574 590614
rect 336954 554614 337574 590058
rect 336954 554058 336986 554614
rect 337542 554058 337574 554614
rect 336954 518614 337574 554058
rect 336954 518058 336986 518614
rect 337542 518058 337574 518614
rect 336954 482614 337574 518058
rect 336954 482058 336986 482614
rect 337542 482058 337574 482614
rect 336954 446614 337574 482058
rect 336954 446058 336986 446614
rect 337542 446058 337574 446614
rect 336954 410614 337574 446058
rect 336954 410058 336986 410614
rect 337542 410058 337574 410614
rect 336954 374614 337574 410058
rect 336954 374058 336986 374614
rect 337542 374058 337574 374614
rect 336954 338614 337574 374058
rect 336954 338058 336986 338614
rect 337542 338058 337574 338614
rect 336954 302614 337574 338058
rect 336954 302058 336986 302614
rect 337542 302058 337574 302614
rect 336954 266614 337574 302058
rect 336954 266058 336986 266614
rect 337542 266058 337574 266614
rect 336954 230614 337574 266058
rect 336954 230058 336986 230614
rect 337542 230058 337574 230614
rect 336954 194614 337574 230058
rect 336954 194058 336986 194614
rect 337542 194058 337574 194614
rect 336954 158614 337574 194058
rect 336954 158058 336986 158614
rect 337542 158058 337574 158614
rect 336954 122614 337574 158058
rect 336954 122058 336986 122614
rect 337542 122058 337574 122614
rect 336954 86614 337574 122058
rect 336954 86058 336986 86614
rect 337542 86058 337574 86614
rect 336954 50614 337574 86058
rect 336954 50058 336986 50614
rect 337542 50058 337574 50614
rect 336954 14614 337574 50058
rect 336954 14058 336986 14614
rect 337542 14058 337574 14614
rect 336954 -3226 337574 14058
rect 336954 -3782 336986 -3226
rect 337542 -3782 337574 -3226
rect 336954 -7654 337574 -3782
rect 340674 708678 341294 711590
rect 340674 708122 340706 708678
rect 341262 708122 341294 708678
rect 340674 666334 341294 708122
rect 340674 665778 340706 666334
rect 341262 665778 341294 666334
rect 340674 630334 341294 665778
rect 340674 629778 340706 630334
rect 341262 629778 341294 630334
rect 340674 594334 341294 629778
rect 340674 593778 340706 594334
rect 341262 593778 341294 594334
rect 340674 558334 341294 593778
rect 340674 557778 340706 558334
rect 341262 557778 341294 558334
rect 340674 522334 341294 557778
rect 340674 521778 340706 522334
rect 341262 521778 341294 522334
rect 340674 486334 341294 521778
rect 340674 485778 340706 486334
rect 341262 485778 341294 486334
rect 340674 450334 341294 485778
rect 340674 449778 340706 450334
rect 341262 449778 341294 450334
rect 340674 414334 341294 449778
rect 340674 413778 340706 414334
rect 341262 413778 341294 414334
rect 340674 378334 341294 413778
rect 340674 377778 340706 378334
rect 341262 377778 341294 378334
rect 340674 342334 341294 377778
rect 340674 341778 340706 342334
rect 341262 341778 341294 342334
rect 340674 306334 341294 341778
rect 340674 305778 340706 306334
rect 341262 305778 341294 306334
rect 340674 270334 341294 305778
rect 340674 269778 340706 270334
rect 341262 269778 341294 270334
rect 340674 234334 341294 269778
rect 340674 233778 340706 234334
rect 341262 233778 341294 234334
rect 340674 198334 341294 233778
rect 340674 197778 340706 198334
rect 341262 197778 341294 198334
rect 340674 162334 341294 197778
rect 340674 161778 340706 162334
rect 341262 161778 341294 162334
rect 340674 126334 341294 161778
rect 340674 125778 340706 126334
rect 341262 125778 341294 126334
rect 340674 90334 341294 125778
rect 340674 89778 340706 90334
rect 341262 89778 341294 90334
rect 340674 54334 341294 89778
rect 340674 53778 340706 54334
rect 341262 53778 341294 54334
rect 340674 18334 341294 53778
rect 340674 17778 340706 18334
rect 341262 17778 341294 18334
rect 340674 -4186 341294 17778
rect 340674 -4742 340706 -4186
rect 341262 -4742 341294 -4186
rect 340674 -7654 341294 -4742
rect 344394 709638 345014 711590
rect 344394 709082 344426 709638
rect 344982 709082 345014 709638
rect 344394 670054 345014 709082
rect 344394 669498 344426 670054
rect 344982 669498 345014 670054
rect 344394 634054 345014 669498
rect 344394 633498 344426 634054
rect 344982 633498 345014 634054
rect 344394 598054 345014 633498
rect 344394 597498 344426 598054
rect 344982 597498 345014 598054
rect 344394 562054 345014 597498
rect 344394 561498 344426 562054
rect 344982 561498 345014 562054
rect 344394 526054 345014 561498
rect 344394 525498 344426 526054
rect 344982 525498 345014 526054
rect 344394 490054 345014 525498
rect 344394 489498 344426 490054
rect 344982 489498 345014 490054
rect 344394 454054 345014 489498
rect 344394 453498 344426 454054
rect 344982 453498 345014 454054
rect 344394 418054 345014 453498
rect 344394 417498 344426 418054
rect 344982 417498 345014 418054
rect 344394 382054 345014 417498
rect 344394 381498 344426 382054
rect 344982 381498 345014 382054
rect 344394 346054 345014 381498
rect 344394 345498 344426 346054
rect 344982 345498 345014 346054
rect 344394 310054 345014 345498
rect 344394 309498 344426 310054
rect 344982 309498 345014 310054
rect 344394 274054 345014 309498
rect 344394 273498 344426 274054
rect 344982 273498 345014 274054
rect 344394 238054 345014 273498
rect 344394 237498 344426 238054
rect 344982 237498 345014 238054
rect 344394 202054 345014 237498
rect 344394 201498 344426 202054
rect 344982 201498 345014 202054
rect 344394 166054 345014 201498
rect 344394 165498 344426 166054
rect 344982 165498 345014 166054
rect 344394 130054 345014 165498
rect 344394 129498 344426 130054
rect 344982 129498 345014 130054
rect 344394 94054 345014 129498
rect 344394 93498 344426 94054
rect 344982 93498 345014 94054
rect 344394 58054 345014 93498
rect 344394 57498 344426 58054
rect 344982 57498 345014 58054
rect 344394 22054 345014 57498
rect 344394 21498 344426 22054
rect 344982 21498 345014 22054
rect 344394 -5146 345014 21498
rect 344394 -5702 344426 -5146
rect 344982 -5702 345014 -5146
rect 344394 -7654 345014 -5702
rect 348114 710598 348734 711590
rect 348114 710042 348146 710598
rect 348702 710042 348734 710598
rect 348114 673774 348734 710042
rect 348114 673218 348146 673774
rect 348702 673218 348734 673774
rect 348114 637774 348734 673218
rect 348114 637218 348146 637774
rect 348702 637218 348734 637774
rect 348114 601774 348734 637218
rect 348114 601218 348146 601774
rect 348702 601218 348734 601774
rect 348114 565774 348734 601218
rect 348114 565218 348146 565774
rect 348702 565218 348734 565774
rect 348114 529774 348734 565218
rect 348114 529218 348146 529774
rect 348702 529218 348734 529774
rect 348114 493774 348734 529218
rect 348114 493218 348146 493774
rect 348702 493218 348734 493774
rect 348114 457774 348734 493218
rect 348114 457218 348146 457774
rect 348702 457218 348734 457774
rect 348114 421774 348734 457218
rect 348114 421218 348146 421774
rect 348702 421218 348734 421774
rect 348114 385774 348734 421218
rect 348114 385218 348146 385774
rect 348702 385218 348734 385774
rect 348114 349774 348734 385218
rect 348114 349218 348146 349774
rect 348702 349218 348734 349774
rect 348114 313774 348734 349218
rect 348114 313218 348146 313774
rect 348702 313218 348734 313774
rect 348114 277774 348734 313218
rect 348114 277218 348146 277774
rect 348702 277218 348734 277774
rect 348114 241774 348734 277218
rect 348114 241218 348146 241774
rect 348702 241218 348734 241774
rect 348114 205774 348734 241218
rect 348114 205218 348146 205774
rect 348702 205218 348734 205774
rect 348114 169774 348734 205218
rect 348114 169218 348146 169774
rect 348702 169218 348734 169774
rect 348114 133774 348734 169218
rect 348114 133218 348146 133774
rect 348702 133218 348734 133774
rect 348114 97774 348734 133218
rect 348114 97218 348146 97774
rect 348702 97218 348734 97774
rect 348114 61774 348734 97218
rect 348114 61218 348146 61774
rect 348702 61218 348734 61774
rect 348114 25774 348734 61218
rect 348114 25218 348146 25774
rect 348702 25218 348734 25774
rect 348114 -6106 348734 25218
rect 348114 -6662 348146 -6106
rect 348702 -6662 348734 -6106
rect 348114 -7654 348734 -6662
rect 351834 711558 352454 711590
rect 351834 711002 351866 711558
rect 352422 711002 352454 711558
rect 351834 677494 352454 711002
rect 351834 676938 351866 677494
rect 352422 676938 352454 677494
rect 351834 641494 352454 676938
rect 351834 640938 351866 641494
rect 352422 640938 352454 641494
rect 351834 605494 352454 640938
rect 351834 604938 351866 605494
rect 352422 604938 352454 605494
rect 351834 569494 352454 604938
rect 351834 568938 351866 569494
rect 352422 568938 352454 569494
rect 351834 533494 352454 568938
rect 351834 532938 351866 533494
rect 352422 532938 352454 533494
rect 351834 497494 352454 532938
rect 351834 496938 351866 497494
rect 352422 496938 352454 497494
rect 351834 461494 352454 496938
rect 351834 460938 351866 461494
rect 352422 460938 352454 461494
rect 351834 425494 352454 460938
rect 351834 424938 351866 425494
rect 352422 424938 352454 425494
rect 351834 389494 352454 424938
rect 351834 388938 351866 389494
rect 352422 388938 352454 389494
rect 351834 353494 352454 388938
rect 351834 352938 351866 353494
rect 352422 352938 352454 353494
rect 351834 317494 352454 352938
rect 351834 316938 351866 317494
rect 352422 316938 352454 317494
rect 351834 281494 352454 316938
rect 351834 280938 351866 281494
rect 352422 280938 352454 281494
rect 351834 245494 352454 280938
rect 351834 244938 351866 245494
rect 352422 244938 352454 245494
rect 351834 209494 352454 244938
rect 351834 208938 351866 209494
rect 352422 208938 352454 209494
rect 351834 173494 352454 208938
rect 351834 172938 351866 173494
rect 352422 172938 352454 173494
rect 351834 137494 352454 172938
rect 351834 136938 351866 137494
rect 352422 136938 352454 137494
rect 351834 101494 352454 136938
rect 351834 100938 351866 101494
rect 352422 100938 352454 101494
rect 351834 65494 352454 100938
rect 351834 64938 351866 65494
rect 352422 64938 352454 65494
rect 351834 29494 352454 64938
rect 351834 28938 351866 29494
rect 352422 28938 352454 29494
rect 351834 -7066 352454 28938
rect 351834 -7622 351866 -7066
rect 352422 -7622 352454 -7066
rect 351834 -7654 352454 -7622
rect 361794 704838 362414 711590
rect 361794 704282 361826 704838
rect 362382 704282 362414 704838
rect 361794 687454 362414 704282
rect 361794 686898 361826 687454
rect 362382 686898 362414 687454
rect 361794 651454 362414 686898
rect 361794 650898 361826 651454
rect 362382 650898 362414 651454
rect 361794 615454 362414 650898
rect 361794 614898 361826 615454
rect 362382 614898 362414 615454
rect 361794 579454 362414 614898
rect 361794 578898 361826 579454
rect 362382 578898 362414 579454
rect 361794 543454 362414 578898
rect 361794 542898 361826 543454
rect 362382 542898 362414 543454
rect 361794 507454 362414 542898
rect 361794 506898 361826 507454
rect 362382 506898 362414 507454
rect 361794 471454 362414 506898
rect 361794 470898 361826 471454
rect 362382 470898 362414 471454
rect 361794 435454 362414 470898
rect 361794 434898 361826 435454
rect 362382 434898 362414 435454
rect 361794 399454 362414 434898
rect 361794 398898 361826 399454
rect 362382 398898 362414 399454
rect 361794 363454 362414 398898
rect 361794 362898 361826 363454
rect 362382 362898 362414 363454
rect 361794 327454 362414 362898
rect 361794 326898 361826 327454
rect 362382 326898 362414 327454
rect 361794 291454 362414 326898
rect 361794 290898 361826 291454
rect 362382 290898 362414 291454
rect 361794 255454 362414 290898
rect 361794 254898 361826 255454
rect 362382 254898 362414 255454
rect 361794 219454 362414 254898
rect 361794 218898 361826 219454
rect 362382 218898 362414 219454
rect 361794 183454 362414 218898
rect 361794 182898 361826 183454
rect 362382 182898 362414 183454
rect 361794 147454 362414 182898
rect 361794 146898 361826 147454
rect 362382 146898 362414 147454
rect 361794 111454 362414 146898
rect 361794 110898 361826 111454
rect 362382 110898 362414 111454
rect 361794 75454 362414 110898
rect 361794 74898 361826 75454
rect 362382 74898 362414 75454
rect 361794 39454 362414 74898
rect 361794 38898 361826 39454
rect 362382 38898 362414 39454
rect 361794 3454 362414 38898
rect 361794 2898 361826 3454
rect 362382 2898 362414 3454
rect 361794 -346 362414 2898
rect 361794 -902 361826 -346
rect 362382 -902 362414 -346
rect 361794 -7654 362414 -902
rect 365514 705798 366134 711590
rect 365514 705242 365546 705798
rect 366102 705242 366134 705798
rect 365514 691174 366134 705242
rect 365514 690618 365546 691174
rect 366102 690618 366134 691174
rect 365514 655174 366134 690618
rect 365514 654618 365546 655174
rect 366102 654618 366134 655174
rect 365514 619174 366134 654618
rect 365514 618618 365546 619174
rect 366102 618618 366134 619174
rect 365514 583174 366134 618618
rect 365514 582618 365546 583174
rect 366102 582618 366134 583174
rect 365514 547174 366134 582618
rect 365514 546618 365546 547174
rect 366102 546618 366134 547174
rect 365514 511174 366134 546618
rect 365514 510618 365546 511174
rect 366102 510618 366134 511174
rect 365514 475174 366134 510618
rect 365514 474618 365546 475174
rect 366102 474618 366134 475174
rect 365514 439174 366134 474618
rect 365514 438618 365546 439174
rect 366102 438618 366134 439174
rect 365514 403174 366134 438618
rect 365514 402618 365546 403174
rect 366102 402618 366134 403174
rect 365514 367174 366134 402618
rect 365514 366618 365546 367174
rect 366102 366618 366134 367174
rect 365514 331174 366134 366618
rect 365514 330618 365546 331174
rect 366102 330618 366134 331174
rect 365514 295174 366134 330618
rect 365514 294618 365546 295174
rect 366102 294618 366134 295174
rect 365514 259174 366134 294618
rect 365514 258618 365546 259174
rect 366102 258618 366134 259174
rect 365514 223174 366134 258618
rect 365514 222618 365546 223174
rect 366102 222618 366134 223174
rect 365514 187174 366134 222618
rect 365514 186618 365546 187174
rect 366102 186618 366134 187174
rect 365514 151174 366134 186618
rect 365514 150618 365546 151174
rect 366102 150618 366134 151174
rect 365514 115174 366134 150618
rect 365514 114618 365546 115174
rect 366102 114618 366134 115174
rect 365514 79174 366134 114618
rect 365514 78618 365546 79174
rect 366102 78618 366134 79174
rect 365514 43174 366134 78618
rect 365514 42618 365546 43174
rect 366102 42618 366134 43174
rect 365514 7174 366134 42618
rect 365514 6618 365546 7174
rect 366102 6618 366134 7174
rect 365514 -1306 366134 6618
rect 365514 -1862 365546 -1306
rect 366102 -1862 366134 -1306
rect 365514 -7654 366134 -1862
rect 369234 706758 369854 711590
rect 369234 706202 369266 706758
rect 369822 706202 369854 706758
rect 369234 694894 369854 706202
rect 369234 694338 369266 694894
rect 369822 694338 369854 694894
rect 369234 658894 369854 694338
rect 369234 658338 369266 658894
rect 369822 658338 369854 658894
rect 369234 622894 369854 658338
rect 369234 622338 369266 622894
rect 369822 622338 369854 622894
rect 369234 586894 369854 622338
rect 369234 586338 369266 586894
rect 369822 586338 369854 586894
rect 369234 550894 369854 586338
rect 369234 550338 369266 550894
rect 369822 550338 369854 550894
rect 369234 514894 369854 550338
rect 369234 514338 369266 514894
rect 369822 514338 369854 514894
rect 369234 478894 369854 514338
rect 369234 478338 369266 478894
rect 369822 478338 369854 478894
rect 369234 442894 369854 478338
rect 369234 442338 369266 442894
rect 369822 442338 369854 442894
rect 369234 406894 369854 442338
rect 369234 406338 369266 406894
rect 369822 406338 369854 406894
rect 369234 370894 369854 406338
rect 369234 370338 369266 370894
rect 369822 370338 369854 370894
rect 369234 334894 369854 370338
rect 369234 334338 369266 334894
rect 369822 334338 369854 334894
rect 369234 298894 369854 334338
rect 369234 298338 369266 298894
rect 369822 298338 369854 298894
rect 369234 262894 369854 298338
rect 369234 262338 369266 262894
rect 369822 262338 369854 262894
rect 369234 226894 369854 262338
rect 369234 226338 369266 226894
rect 369822 226338 369854 226894
rect 369234 190894 369854 226338
rect 369234 190338 369266 190894
rect 369822 190338 369854 190894
rect 369234 154894 369854 190338
rect 369234 154338 369266 154894
rect 369822 154338 369854 154894
rect 369234 118894 369854 154338
rect 369234 118338 369266 118894
rect 369822 118338 369854 118894
rect 369234 82894 369854 118338
rect 369234 82338 369266 82894
rect 369822 82338 369854 82894
rect 369234 46894 369854 82338
rect 369234 46338 369266 46894
rect 369822 46338 369854 46894
rect 369234 10894 369854 46338
rect 369234 10338 369266 10894
rect 369822 10338 369854 10894
rect 369234 -2266 369854 10338
rect 369234 -2822 369266 -2266
rect 369822 -2822 369854 -2266
rect 369234 -7654 369854 -2822
rect 372954 707718 373574 711590
rect 372954 707162 372986 707718
rect 373542 707162 373574 707718
rect 372954 698614 373574 707162
rect 372954 698058 372986 698614
rect 373542 698058 373574 698614
rect 372954 662614 373574 698058
rect 372954 662058 372986 662614
rect 373542 662058 373574 662614
rect 372954 626614 373574 662058
rect 372954 626058 372986 626614
rect 373542 626058 373574 626614
rect 372954 590614 373574 626058
rect 372954 590058 372986 590614
rect 373542 590058 373574 590614
rect 372954 554614 373574 590058
rect 372954 554058 372986 554614
rect 373542 554058 373574 554614
rect 372954 518614 373574 554058
rect 372954 518058 372986 518614
rect 373542 518058 373574 518614
rect 372954 482614 373574 518058
rect 372954 482058 372986 482614
rect 373542 482058 373574 482614
rect 372954 446614 373574 482058
rect 372954 446058 372986 446614
rect 373542 446058 373574 446614
rect 372954 410614 373574 446058
rect 372954 410058 372986 410614
rect 373542 410058 373574 410614
rect 372954 374614 373574 410058
rect 372954 374058 372986 374614
rect 373542 374058 373574 374614
rect 372954 338614 373574 374058
rect 372954 338058 372986 338614
rect 373542 338058 373574 338614
rect 372954 302614 373574 338058
rect 372954 302058 372986 302614
rect 373542 302058 373574 302614
rect 372954 266614 373574 302058
rect 372954 266058 372986 266614
rect 373542 266058 373574 266614
rect 372954 230614 373574 266058
rect 372954 230058 372986 230614
rect 373542 230058 373574 230614
rect 372954 194614 373574 230058
rect 372954 194058 372986 194614
rect 373542 194058 373574 194614
rect 372954 158614 373574 194058
rect 372954 158058 372986 158614
rect 373542 158058 373574 158614
rect 372954 122614 373574 158058
rect 372954 122058 372986 122614
rect 373542 122058 373574 122614
rect 372954 86614 373574 122058
rect 372954 86058 372986 86614
rect 373542 86058 373574 86614
rect 372954 50614 373574 86058
rect 372954 50058 372986 50614
rect 373542 50058 373574 50614
rect 372954 14614 373574 50058
rect 372954 14058 372986 14614
rect 373542 14058 373574 14614
rect 372954 -3226 373574 14058
rect 372954 -3782 372986 -3226
rect 373542 -3782 373574 -3226
rect 372954 -7654 373574 -3782
rect 376674 708678 377294 711590
rect 376674 708122 376706 708678
rect 377262 708122 377294 708678
rect 376674 666334 377294 708122
rect 376674 665778 376706 666334
rect 377262 665778 377294 666334
rect 376674 630334 377294 665778
rect 376674 629778 376706 630334
rect 377262 629778 377294 630334
rect 376674 594334 377294 629778
rect 376674 593778 376706 594334
rect 377262 593778 377294 594334
rect 376674 558334 377294 593778
rect 376674 557778 376706 558334
rect 377262 557778 377294 558334
rect 376674 522334 377294 557778
rect 376674 521778 376706 522334
rect 377262 521778 377294 522334
rect 376674 486334 377294 521778
rect 376674 485778 376706 486334
rect 377262 485778 377294 486334
rect 376674 450334 377294 485778
rect 376674 449778 376706 450334
rect 377262 449778 377294 450334
rect 376674 414334 377294 449778
rect 376674 413778 376706 414334
rect 377262 413778 377294 414334
rect 376674 378334 377294 413778
rect 376674 377778 376706 378334
rect 377262 377778 377294 378334
rect 376674 342334 377294 377778
rect 376674 341778 376706 342334
rect 377262 341778 377294 342334
rect 376674 306334 377294 341778
rect 376674 305778 376706 306334
rect 377262 305778 377294 306334
rect 376674 270334 377294 305778
rect 376674 269778 376706 270334
rect 377262 269778 377294 270334
rect 376674 234334 377294 269778
rect 376674 233778 376706 234334
rect 377262 233778 377294 234334
rect 376674 198334 377294 233778
rect 376674 197778 376706 198334
rect 377262 197778 377294 198334
rect 376674 162334 377294 197778
rect 376674 161778 376706 162334
rect 377262 161778 377294 162334
rect 376674 126334 377294 161778
rect 376674 125778 376706 126334
rect 377262 125778 377294 126334
rect 376674 90334 377294 125778
rect 376674 89778 376706 90334
rect 377262 89778 377294 90334
rect 376674 54334 377294 89778
rect 376674 53778 376706 54334
rect 377262 53778 377294 54334
rect 376674 18334 377294 53778
rect 376674 17778 376706 18334
rect 377262 17778 377294 18334
rect 376674 -4186 377294 17778
rect 376674 -4742 376706 -4186
rect 377262 -4742 377294 -4186
rect 376674 -7654 377294 -4742
rect 380394 709638 381014 711590
rect 380394 709082 380426 709638
rect 380982 709082 381014 709638
rect 380394 670054 381014 709082
rect 380394 669498 380426 670054
rect 380982 669498 381014 670054
rect 380394 634054 381014 669498
rect 380394 633498 380426 634054
rect 380982 633498 381014 634054
rect 380394 598054 381014 633498
rect 380394 597498 380426 598054
rect 380982 597498 381014 598054
rect 380394 562054 381014 597498
rect 380394 561498 380426 562054
rect 380982 561498 381014 562054
rect 380394 526054 381014 561498
rect 380394 525498 380426 526054
rect 380982 525498 381014 526054
rect 380394 490054 381014 525498
rect 380394 489498 380426 490054
rect 380982 489498 381014 490054
rect 380394 454054 381014 489498
rect 380394 453498 380426 454054
rect 380982 453498 381014 454054
rect 380394 418054 381014 453498
rect 380394 417498 380426 418054
rect 380982 417498 381014 418054
rect 380394 382054 381014 417498
rect 380394 381498 380426 382054
rect 380982 381498 381014 382054
rect 380394 346054 381014 381498
rect 380394 345498 380426 346054
rect 380982 345498 381014 346054
rect 380394 310054 381014 345498
rect 380394 309498 380426 310054
rect 380982 309498 381014 310054
rect 380394 274054 381014 309498
rect 380394 273498 380426 274054
rect 380982 273498 381014 274054
rect 380394 238054 381014 273498
rect 380394 237498 380426 238054
rect 380982 237498 381014 238054
rect 380394 202054 381014 237498
rect 380394 201498 380426 202054
rect 380982 201498 381014 202054
rect 380394 166054 381014 201498
rect 380394 165498 380426 166054
rect 380982 165498 381014 166054
rect 380394 130054 381014 165498
rect 380394 129498 380426 130054
rect 380982 129498 381014 130054
rect 380394 94054 381014 129498
rect 380394 93498 380426 94054
rect 380982 93498 381014 94054
rect 380394 58054 381014 93498
rect 380394 57498 380426 58054
rect 380982 57498 381014 58054
rect 380394 22054 381014 57498
rect 380394 21498 380426 22054
rect 380982 21498 381014 22054
rect 380394 -5146 381014 21498
rect 380394 -5702 380426 -5146
rect 380982 -5702 381014 -5146
rect 380394 -7654 381014 -5702
rect 384114 710598 384734 711590
rect 384114 710042 384146 710598
rect 384702 710042 384734 710598
rect 384114 673774 384734 710042
rect 384114 673218 384146 673774
rect 384702 673218 384734 673774
rect 384114 637774 384734 673218
rect 384114 637218 384146 637774
rect 384702 637218 384734 637774
rect 384114 601774 384734 637218
rect 384114 601218 384146 601774
rect 384702 601218 384734 601774
rect 384114 565774 384734 601218
rect 384114 565218 384146 565774
rect 384702 565218 384734 565774
rect 384114 529774 384734 565218
rect 384114 529218 384146 529774
rect 384702 529218 384734 529774
rect 384114 493774 384734 529218
rect 384114 493218 384146 493774
rect 384702 493218 384734 493774
rect 384114 457774 384734 493218
rect 384114 457218 384146 457774
rect 384702 457218 384734 457774
rect 384114 421774 384734 457218
rect 384114 421218 384146 421774
rect 384702 421218 384734 421774
rect 384114 385774 384734 421218
rect 384114 385218 384146 385774
rect 384702 385218 384734 385774
rect 384114 349774 384734 385218
rect 384114 349218 384146 349774
rect 384702 349218 384734 349774
rect 384114 313774 384734 349218
rect 384114 313218 384146 313774
rect 384702 313218 384734 313774
rect 384114 277774 384734 313218
rect 384114 277218 384146 277774
rect 384702 277218 384734 277774
rect 384114 241774 384734 277218
rect 384114 241218 384146 241774
rect 384702 241218 384734 241774
rect 384114 205774 384734 241218
rect 384114 205218 384146 205774
rect 384702 205218 384734 205774
rect 384114 169774 384734 205218
rect 384114 169218 384146 169774
rect 384702 169218 384734 169774
rect 384114 133774 384734 169218
rect 384114 133218 384146 133774
rect 384702 133218 384734 133774
rect 384114 97774 384734 133218
rect 384114 97218 384146 97774
rect 384702 97218 384734 97774
rect 384114 61774 384734 97218
rect 384114 61218 384146 61774
rect 384702 61218 384734 61774
rect 384114 25774 384734 61218
rect 384114 25218 384146 25774
rect 384702 25218 384734 25774
rect 384114 -6106 384734 25218
rect 384114 -6662 384146 -6106
rect 384702 -6662 384734 -6106
rect 384114 -7654 384734 -6662
rect 387834 711558 388454 711590
rect 387834 711002 387866 711558
rect 388422 711002 388454 711558
rect 387834 677494 388454 711002
rect 387834 676938 387866 677494
rect 388422 676938 388454 677494
rect 387834 641494 388454 676938
rect 387834 640938 387866 641494
rect 388422 640938 388454 641494
rect 387834 605494 388454 640938
rect 387834 604938 387866 605494
rect 388422 604938 388454 605494
rect 387834 569494 388454 604938
rect 387834 568938 387866 569494
rect 388422 568938 388454 569494
rect 387834 533494 388454 568938
rect 387834 532938 387866 533494
rect 388422 532938 388454 533494
rect 387834 497494 388454 532938
rect 387834 496938 387866 497494
rect 388422 496938 388454 497494
rect 387834 461494 388454 496938
rect 387834 460938 387866 461494
rect 388422 460938 388454 461494
rect 387834 425494 388454 460938
rect 387834 424938 387866 425494
rect 388422 424938 388454 425494
rect 387834 389494 388454 424938
rect 387834 388938 387866 389494
rect 388422 388938 388454 389494
rect 387834 353494 388454 388938
rect 387834 352938 387866 353494
rect 388422 352938 388454 353494
rect 387834 317494 388454 352938
rect 387834 316938 387866 317494
rect 388422 316938 388454 317494
rect 387834 281494 388454 316938
rect 387834 280938 387866 281494
rect 388422 280938 388454 281494
rect 387834 245494 388454 280938
rect 387834 244938 387866 245494
rect 388422 244938 388454 245494
rect 387834 209494 388454 244938
rect 387834 208938 387866 209494
rect 388422 208938 388454 209494
rect 387834 173494 388454 208938
rect 387834 172938 387866 173494
rect 388422 172938 388454 173494
rect 387834 137494 388454 172938
rect 387834 136938 387866 137494
rect 388422 136938 388454 137494
rect 387834 101494 388454 136938
rect 387834 100938 387866 101494
rect 388422 100938 388454 101494
rect 387834 65494 388454 100938
rect 387834 64938 387866 65494
rect 388422 64938 388454 65494
rect 387834 29494 388454 64938
rect 387834 28938 387866 29494
rect 388422 28938 388454 29494
rect 387834 -7066 388454 28938
rect 387834 -7622 387866 -7066
rect 388422 -7622 388454 -7066
rect 387834 -7654 388454 -7622
rect 397794 704838 398414 711590
rect 397794 704282 397826 704838
rect 398382 704282 398414 704838
rect 397794 687454 398414 704282
rect 397794 686898 397826 687454
rect 398382 686898 398414 687454
rect 397794 651454 398414 686898
rect 397794 650898 397826 651454
rect 398382 650898 398414 651454
rect 397794 615454 398414 650898
rect 397794 614898 397826 615454
rect 398382 614898 398414 615454
rect 397794 579454 398414 614898
rect 397794 578898 397826 579454
rect 398382 578898 398414 579454
rect 397794 543454 398414 578898
rect 397794 542898 397826 543454
rect 398382 542898 398414 543454
rect 397794 507454 398414 542898
rect 397794 506898 397826 507454
rect 398382 506898 398414 507454
rect 397794 471454 398414 506898
rect 397794 470898 397826 471454
rect 398382 470898 398414 471454
rect 397794 435454 398414 470898
rect 397794 434898 397826 435454
rect 398382 434898 398414 435454
rect 397794 399454 398414 434898
rect 397794 398898 397826 399454
rect 398382 398898 398414 399454
rect 397794 363454 398414 398898
rect 397794 362898 397826 363454
rect 398382 362898 398414 363454
rect 397794 327454 398414 362898
rect 397794 326898 397826 327454
rect 398382 326898 398414 327454
rect 397794 291454 398414 326898
rect 397794 290898 397826 291454
rect 398382 290898 398414 291454
rect 397794 255454 398414 290898
rect 397794 254898 397826 255454
rect 398382 254898 398414 255454
rect 397794 219454 398414 254898
rect 397794 218898 397826 219454
rect 398382 218898 398414 219454
rect 397794 183454 398414 218898
rect 397794 182898 397826 183454
rect 398382 182898 398414 183454
rect 397794 147454 398414 182898
rect 397794 146898 397826 147454
rect 398382 146898 398414 147454
rect 397794 111454 398414 146898
rect 397794 110898 397826 111454
rect 398382 110898 398414 111454
rect 397794 75454 398414 110898
rect 397794 74898 397826 75454
rect 398382 74898 398414 75454
rect 397794 39454 398414 74898
rect 397794 38898 397826 39454
rect 398382 38898 398414 39454
rect 397794 3454 398414 38898
rect 397794 2898 397826 3454
rect 398382 2898 398414 3454
rect 397794 -346 398414 2898
rect 397794 -902 397826 -346
rect 398382 -902 398414 -346
rect 397794 -7654 398414 -902
rect 401514 705798 402134 711590
rect 401514 705242 401546 705798
rect 402102 705242 402134 705798
rect 401514 691174 402134 705242
rect 401514 690618 401546 691174
rect 402102 690618 402134 691174
rect 401514 655174 402134 690618
rect 401514 654618 401546 655174
rect 402102 654618 402134 655174
rect 401514 619174 402134 654618
rect 401514 618618 401546 619174
rect 402102 618618 402134 619174
rect 401514 583174 402134 618618
rect 401514 582618 401546 583174
rect 402102 582618 402134 583174
rect 401514 547174 402134 582618
rect 401514 546618 401546 547174
rect 402102 546618 402134 547174
rect 401514 511174 402134 546618
rect 401514 510618 401546 511174
rect 402102 510618 402134 511174
rect 401514 475174 402134 510618
rect 401514 474618 401546 475174
rect 402102 474618 402134 475174
rect 401514 439174 402134 474618
rect 401514 438618 401546 439174
rect 402102 438618 402134 439174
rect 401514 403174 402134 438618
rect 401514 402618 401546 403174
rect 402102 402618 402134 403174
rect 401514 367174 402134 402618
rect 401514 366618 401546 367174
rect 402102 366618 402134 367174
rect 401514 331174 402134 366618
rect 401514 330618 401546 331174
rect 402102 330618 402134 331174
rect 401514 295174 402134 330618
rect 401514 294618 401546 295174
rect 402102 294618 402134 295174
rect 401514 259174 402134 294618
rect 401514 258618 401546 259174
rect 402102 258618 402134 259174
rect 401514 223174 402134 258618
rect 401514 222618 401546 223174
rect 402102 222618 402134 223174
rect 401514 187174 402134 222618
rect 401514 186618 401546 187174
rect 402102 186618 402134 187174
rect 401514 151174 402134 186618
rect 401514 150618 401546 151174
rect 402102 150618 402134 151174
rect 401514 115174 402134 150618
rect 401514 114618 401546 115174
rect 402102 114618 402134 115174
rect 401514 79174 402134 114618
rect 401514 78618 401546 79174
rect 402102 78618 402134 79174
rect 401514 43174 402134 78618
rect 401514 42618 401546 43174
rect 402102 42618 402134 43174
rect 401514 7174 402134 42618
rect 401514 6618 401546 7174
rect 402102 6618 402134 7174
rect 401514 -1306 402134 6618
rect 401514 -1862 401546 -1306
rect 402102 -1862 402134 -1306
rect 401514 -7654 402134 -1862
rect 405234 706758 405854 711590
rect 405234 706202 405266 706758
rect 405822 706202 405854 706758
rect 405234 694894 405854 706202
rect 405234 694338 405266 694894
rect 405822 694338 405854 694894
rect 405234 658894 405854 694338
rect 405234 658338 405266 658894
rect 405822 658338 405854 658894
rect 405234 622894 405854 658338
rect 405234 622338 405266 622894
rect 405822 622338 405854 622894
rect 405234 586894 405854 622338
rect 405234 586338 405266 586894
rect 405822 586338 405854 586894
rect 405234 550894 405854 586338
rect 405234 550338 405266 550894
rect 405822 550338 405854 550894
rect 405234 514894 405854 550338
rect 405234 514338 405266 514894
rect 405822 514338 405854 514894
rect 405234 478894 405854 514338
rect 405234 478338 405266 478894
rect 405822 478338 405854 478894
rect 405234 442894 405854 478338
rect 405234 442338 405266 442894
rect 405822 442338 405854 442894
rect 405234 406894 405854 442338
rect 405234 406338 405266 406894
rect 405822 406338 405854 406894
rect 405234 370894 405854 406338
rect 405234 370338 405266 370894
rect 405822 370338 405854 370894
rect 405234 334894 405854 370338
rect 405234 334338 405266 334894
rect 405822 334338 405854 334894
rect 405234 298894 405854 334338
rect 405234 298338 405266 298894
rect 405822 298338 405854 298894
rect 405234 262894 405854 298338
rect 405234 262338 405266 262894
rect 405822 262338 405854 262894
rect 405234 226894 405854 262338
rect 405234 226338 405266 226894
rect 405822 226338 405854 226894
rect 405234 190894 405854 226338
rect 405234 190338 405266 190894
rect 405822 190338 405854 190894
rect 405234 154894 405854 190338
rect 405234 154338 405266 154894
rect 405822 154338 405854 154894
rect 405234 118894 405854 154338
rect 405234 118338 405266 118894
rect 405822 118338 405854 118894
rect 405234 82894 405854 118338
rect 405234 82338 405266 82894
rect 405822 82338 405854 82894
rect 405234 46894 405854 82338
rect 405234 46338 405266 46894
rect 405822 46338 405854 46894
rect 405234 10894 405854 46338
rect 405234 10338 405266 10894
rect 405822 10338 405854 10894
rect 405234 -2266 405854 10338
rect 405234 -2822 405266 -2266
rect 405822 -2822 405854 -2266
rect 405234 -7654 405854 -2822
rect 408954 707718 409574 711590
rect 408954 707162 408986 707718
rect 409542 707162 409574 707718
rect 408954 698614 409574 707162
rect 408954 698058 408986 698614
rect 409542 698058 409574 698614
rect 408954 662614 409574 698058
rect 408954 662058 408986 662614
rect 409542 662058 409574 662614
rect 408954 626614 409574 662058
rect 408954 626058 408986 626614
rect 409542 626058 409574 626614
rect 408954 590614 409574 626058
rect 408954 590058 408986 590614
rect 409542 590058 409574 590614
rect 408954 554614 409574 590058
rect 408954 554058 408986 554614
rect 409542 554058 409574 554614
rect 408954 518614 409574 554058
rect 408954 518058 408986 518614
rect 409542 518058 409574 518614
rect 408954 482614 409574 518058
rect 408954 482058 408986 482614
rect 409542 482058 409574 482614
rect 408954 446614 409574 482058
rect 408954 446058 408986 446614
rect 409542 446058 409574 446614
rect 408954 410614 409574 446058
rect 408954 410058 408986 410614
rect 409542 410058 409574 410614
rect 408954 374614 409574 410058
rect 408954 374058 408986 374614
rect 409542 374058 409574 374614
rect 408954 338614 409574 374058
rect 408954 338058 408986 338614
rect 409542 338058 409574 338614
rect 408954 302614 409574 338058
rect 408954 302058 408986 302614
rect 409542 302058 409574 302614
rect 408954 266614 409574 302058
rect 408954 266058 408986 266614
rect 409542 266058 409574 266614
rect 408954 230614 409574 266058
rect 408954 230058 408986 230614
rect 409542 230058 409574 230614
rect 408954 194614 409574 230058
rect 408954 194058 408986 194614
rect 409542 194058 409574 194614
rect 408954 158614 409574 194058
rect 408954 158058 408986 158614
rect 409542 158058 409574 158614
rect 408954 122614 409574 158058
rect 408954 122058 408986 122614
rect 409542 122058 409574 122614
rect 408954 86614 409574 122058
rect 408954 86058 408986 86614
rect 409542 86058 409574 86614
rect 408954 50614 409574 86058
rect 408954 50058 408986 50614
rect 409542 50058 409574 50614
rect 408954 14614 409574 50058
rect 408954 14058 408986 14614
rect 409542 14058 409574 14614
rect 408954 -3226 409574 14058
rect 408954 -3782 408986 -3226
rect 409542 -3782 409574 -3226
rect 408954 -7654 409574 -3782
rect 412674 708678 413294 711590
rect 412674 708122 412706 708678
rect 413262 708122 413294 708678
rect 412674 666334 413294 708122
rect 412674 665778 412706 666334
rect 413262 665778 413294 666334
rect 412674 630334 413294 665778
rect 412674 629778 412706 630334
rect 413262 629778 413294 630334
rect 412674 594334 413294 629778
rect 412674 593778 412706 594334
rect 413262 593778 413294 594334
rect 412674 558334 413294 593778
rect 412674 557778 412706 558334
rect 413262 557778 413294 558334
rect 412674 522334 413294 557778
rect 412674 521778 412706 522334
rect 413262 521778 413294 522334
rect 412674 486334 413294 521778
rect 412674 485778 412706 486334
rect 413262 485778 413294 486334
rect 412674 450334 413294 485778
rect 412674 449778 412706 450334
rect 413262 449778 413294 450334
rect 412674 414334 413294 449778
rect 412674 413778 412706 414334
rect 413262 413778 413294 414334
rect 412674 378334 413294 413778
rect 412674 377778 412706 378334
rect 413262 377778 413294 378334
rect 412674 342334 413294 377778
rect 412674 341778 412706 342334
rect 413262 341778 413294 342334
rect 412674 306334 413294 341778
rect 412674 305778 412706 306334
rect 413262 305778 413294 306334
rect 412674 270334 413294 305778
rect 412674 269778 412706 270334
rect 413262 269778 413294 270334
rect 412674 234334 413294 269778
rect 412674 233778 412706 234334
rect 413262 233778 413294 234334
rect 412674 198334 413294 233778
rect 412674 197778 412706 198334
rect 413262 197778 413294 198334
rect 412674 162334 413294 197778
rect 412674 161778 412706 162334
rect 413262 161778 413294 162334
rect 412674 126334 413294 161778
rect 412674 125778 412706 126334
rect 413262 125778 413294 126334
rect 412674 90334 413294 125778
rect 412674 89778 412706 90334
rect 413262 89778 413294 90334
rect 412674 54334 413294 89778
rect 412674 53778 412706 54334
rect 413262 53778 413294 54334
rect 412674 18334 413294 53778
rect 412674 17778 412706 18334
rect 413262 17778 413294 18334
rect 412674 -4186 413294 17778
rect 412674 -4742 412706 -4186
rect 413262 -4742 413294 -4186
rect 412674 -7654 413294 -4742
rect 416394 709638 417014 711590
rect 416394 709082 416426 709638
rect 416982 709082 417014 709638
rect 416394 670054 417014 709082
rect 416394 669498 416426 670054
rect 416982 669498 417014 670054
rect 416394 634054 417014 669498
rect 416394 633498 416426 634054
rect 416982 633498 417014 634054
rect 416394 598054 417014 633498
rect 416394 597498 416426 598054
rect 416982 597498 417014 598054
rect 416394 562054 417014 597498
rect 416394 561498 416426 562054
rect 416982 561498 417014 562054
rect 416394 526054 417014 561498
rect 416394 525498 416426 526054
rect 416982 525498 417014 526054
rect 416394 490054 417014 525498
rect 416394 489498 416426 490054
rect 416982 489498 417014 490054
rect 416394 454054 417014 489498
rect 416394 453498 416426 454054
rect 416982 453498 417014 454054
rect 416394 418054 417014 453498
rect 416394 417498 416426 418054
rect 416982 417498 417014 418054
rect 416394 382054 417014 417498
rect 416394 381498 416426 382054
rect 416982 381498 417014 382054
rect 416394 346054 417014 381498
rect 416394 345498 416426 346054
rect 416982 345498 417014 346054
rect 416394 310054 417014 345498
rect 416394 309498 416426 310054
rect 416982 309498 417014 310054
rect 416394 274054 417014 309498
rect 416394 273498 416426 274054
rect 416982 273498 417014 274054
rect 416394 238054 417014 273498
rect 416394 237498 416426 238054
rect 416982 237498 417014 238054
rect 416394 202054 417014 237498
rect 416394 201498 416426 202054
rect 416982 201498 417014 202054
rect 416394 166054 417014 201498
rect 416394 165498 416426 166054
rect 416982 165498 417014 166054
rect 416394 130054 417014 165498
rect 416394 129498 416426 130054
rect 416982 129498 417014 130054
rect 416394 94054 417014 129498
rect 416394 93498 416426 94054
rect 416982 93498 417014 94054
rect 416394 58054 417014 93498
rect 416394 57498 416426 58054
rect 416982 57498 417014 58054
rect 416394 22054 417014 57498
rect 416394 21498 416426 22054
rect 416982 21498 417014 22054
rect 416394 -5146 417014 21498
rect 416394 -5702 416426 -5146
rect 416982 -5702 417014 -5146
rect 416394 -7654 417014 -5702
rect 420114 710598 420734 711590
rect 420114 710042 420146 710598
rect 420702 710042 420734 710598
rect 420114 673774 420734 710042
rect 420114 673218 420146 673774
rect 420702 673218 420734 673774
rect 420114 637774 420734 673218
rect 420114 637218 420146 637774
rect 420702 637218 420734 637774
rect 420114 601774 420734 637218
rect 420114 601218 420146 601774
rect 420702 601218 420734 601774
rect 420114 565774 420734 601218
rect 420114 565218 420146 565774
rect 420702 565218 420734 565774
rect 420114 529774 420734 565218
rect 420114 529218 420146 529774
rect 420702 529218 420734 529774
rect 420114 493774 420734 529218
rect 420114 493218 420146 493774
rect 420702 493218 420734 493774
rect 420114 457774 420734 493218
rect 420114 457218 420146 457774
rect 420702 457218 420734 457774
rect 420114 421774 420734 457218
rect 420114 421218 420146 421774
rect 420702 421218 420734 421774
rect 420114 385774 420734 421218
rect 420114 385218 420146 385774
rect 420702 385218 420734 385774
rect 420114 349774 420734 385218
rect 420114 349218 420146 349774
rect 420702 349218 420734 349774
rect 420114 313774 420734 349218
rect 420114 313218 420146 313774
rect 420702 313218 420734 313774
rect 420114 277774 420734 313218
rect 420114 277218 420146 277774
rect 420702 277218 420734 277774
rect 420114 241774 420734 277218
rect 420114 241218 420146 241774
rect 420702 241218 420734 241774
rect 420114 205774 420734 241218
rect 420114 205218 420146 205774
rect 420702 205218 420734 205774
rect 420114 169774 420734 205218
rect 420114 169218 420146 169774
rect 420702 169218 420734 169774
rect 420114 133774 420734 169218
rect 420114 133218 420146 133774
rect 420702 133218 420734 133774
rect 420114 97774 420734 133218
rect 420114 97218 420146 97774
rect 420702 97218 420734 97774
rect 420114 61774 420734 97218
rect 420114 61218 420146 61774
rect 420702 61218 420734 61774
rect 420114 25774 420734 61218
rect 420114 25218 420146 25774
rect 420702 25218 420734 25774
rect 420114 -6106 420734 25218
rect 420114 -6662 420146 -6106
rect 420702 -6662 420734 -6106
rect 420114 -7654 420734 -6662
rect 423834 711558 424454 711590
rect 423834 711002 423866 711558
rect 424422 711002 424454 711558
rect 423834 677494 424454 711002
rect 423834 676938 423866 677494
rect 424422 676938 424454 677494
rect 423834 641494 424454 676938
rect 423834 640938 423866 641494
rect 424422 640938 424454 641494
rect 423834 605494 424454 640938
rect 423834 604938 423866 605494
rect 424422 604938 424454 605494
rect 423834 569494 424454 604938
rect 423834 568938 423866 569494
rect 424422 568938 424454 569494
rect 423834 533494 424454 568938
rect 423834 532938 423866 533494
rect 424422 532938 424454 533494
rect 423834 497494 424454 532938
rect 423834 496938 423866 497494
rect 424422 496938 424454 497494
rect 423834 461494 424454 496938
rect 423834 460938 423866 461494
rect 424422 460938 424454 461494
rect 423834 425494 424454 460938
rect 423834 424938 423866 425494
rect 424422 424938 424454 425494
rect 423834 389494 424454 424938
rect 423834 388938 423866 389494
rect 424422 388938 424454 389494
rect 423834 353494 424454 388938
rect 423834 352938 423866 353494
rect 424422 352938 424454 353494
rect 423834 317494 424454 352938
rect 423834 316938 423866 317494
rect 424422 316938 424454 317494
rect 423834 281494 424454 316938
rect 423834 280938 423866 281494
rect 424422 280938 424454 281494
rect 423834 245494 424454 280938
rect 423834 244938 423866 245494
rect 424422 244938 424454 245494
rect 423834 209494 424454 244938
rect 423834 208938 423866 209494
rect 424422 208938 424454 209494
rect 423834 173494 424454 208938
rect 423834 172938 423866 173494
rect 424422 172938 424454 173494
rect 423834 137494 424454 172938
rect 423834 136938 423866 137494
rect 424422 136938 424454 137494
rect 423834 101494 424454 136938
rect 423834 100938 423866 101494
rect 424422 100938 424454 101494
rect 423834 65494 424454 100938
rect 423834 64938 423866 65494
rect 424422 64938 424454 65494
rect 423834 29494 424454 64938
rect 423834 28938 423866 29494
rect 424422 28938 424454 29494
rect 423834 -7066 424454 28938
rect 423834 -7622 423866 -7066
rect 424422 -7622 424454 -7066
rect 423834 -7654 424454 -7622
rect 433794 704838 434414 711590
rect 433794 704282 433826 704838
rect 434382 704282 434414 704838
rect 433794 687454 434414 704282
rect 433794 686898 433826 687454
rect 434382 686898 434414 687454
rect 433794 651454 434414 686898
rect 433794 650898 433826 651454
rect 434382 650898 434414 651454
rect 433794 615454 434414 650898
rect 433794 614898 433826 615454
rect 434382 614898 434414 615454
rect 433794 579454 434414 614898
rect 433794 578898 433826 579454
rect 434382 578898 434414 579454
rect 433794 543454 434414 578898
rect 433794 542898 433826 543454
rect 434382 542898 434414 543454
rect 433794 507454 434414 542898
rect 433794 506898 433826 507454
rect 434382 506898 434414 507454
rect 433794 471454 434414 506898
rect 433794 470898 433826 471454
rect 434382 470898 434414 471454
rect 433794 435454 434414 470898
rect 433794 434898 433826 435454
rect 434382 434898 434414 435454
rect 433794 399454 434414 434898
rect 433794 398898 433826 399454
rect 434382 398898 434414 399454
rect 433794 363454 434414 398898
rect 433794 362898 433826 363454
rect 434382 362898 434414 363454
rect 433794 327454 434414 362898
rect 433794 326898 433826 327454
rect 434382 326898 434414 327454
rect 433794 291454 434414 326898
rect 433794 290898 433826 291454
rect 434382 290898 434414 291454
rect 433794 255454 434414 290898
rect 433794 254898 433826 255454
rect 434382 254898 434414 255454
rect 433794 219454 434414 254898
rect 433794 218898 433826 219454
rect 434382 218898 434414 219454
rect 433794 183454 434414 218898
rect 433794 182898 433826 183454
rect 434382 182898 434414 183454
rect 433794 147454 434414 182898
rect 433794 146898 433826 147454
rect 434382 146898 434414 147454
rect 433794 111454 434414 146898
rect 433794 110898 433826 111454
rect 434382 110898 434414 111454
rect 433794 75454 434414 110898
rect 433794 74898 433826 75454
rect 434382 74898 434414 75454
rect 433794 39454 434414 74898
rect 433794 38898 433826 39454
rect 434382 38898 434414 39454
rect 433794 3454 434414 38898
rect 433794 2898 433826 3454
rect 434382 2898 434414 3454
rect 433794 -346 434414 2898
rect 433794 -902 433826 -346
rect 434382 -902 434414 -346
rect 433794 -7654 434414 -902
rect 437514 705798 438134 711590
rect 437514 705242 437546 705798
rect 438102 705242 438134 705798
rect 437514 691174 438134 705242
rect 437514 690618 437546 691174
rect 438102 690618 438134 691174
rect 437514 655174 438134 690618
rect 437514 654618 437546 655174
rect 438102 654618 438134 655174
rect 437514 619174 438134 654618
rect 437514 618618 437546 619174
rect 438102 618618 438134 619174
rect 437514 583174 438134 618618
rect 437514 582618 437546 583174
rect 438102 582618 438134 583174
rect 437514 547174 438134 582618
rect 437514 546618 437546 547174
rect 438102 546618 438134 547174
rect 437514 511174 438134 546618
rect 437514 510618 437546 511174
rect 438102 510618 438134 511174
rect 437514 475174 438134 510618
rect 437514 474618 437546 475174
rect 438102 474618 438134 475174
rect 437514 439174 438134 474618
rect 437514 438618 437546 439174
rect 438102 438618 438134 439174
rect 437514 403174 438134 438618
rect 437514 402618 437546 403174
rect 438102 402618 438134 403174
rect 437514 367174 438134 402618
rect 437514 366618 437546 367174
rect 438102 366618 438134 367174
rect 437514 331174 438134 366618
rect 437514 330618 437546 331174
rect 438102 330618 438134 331174
rect 437514 295174 438134 330618
rect 437514 294618 437546 295174
rect 438102 294618 438134 295174
rect 437514 259174 438134 294618
rect 437514 258618 437546 259174
rect 438102 258618 438134 259174
rect 437514 223174 438134 258618
rect 437514 222618 437546 223174
rect 438102 222618 438134 223174
rect 437514 187174 438134 222618
rect 437514 186618 437546 187174
rect 438102 186618 438134 187174
rect 437514 151174 438134 186618
rect 437514 150618 437546 151174
rect 438102 150618 438134 151174
rect 437514 115174 438134 150618
rect 437514 114618 437546 115174
rect 438102 114618 438134 115174
rect 437514 79174 438134 114618
rect 437514 78618 437546 79174
rect 438102 78618 438134 79174
rect 437514 43174 438134 78618
rect 437514 42618 437546 43174
rect 438102 42618 438134 43174
rect 437514 7174 438134 42618
rect 437514 6618 437546 7174
rect 438102 6618 438134 7174
rect 437514 -1306 438134 6618
rect 437514 -1862 437546 -1306
rect 438102 -1862 438134 -1306
rect 437514 -7654 438134 -1862
rect 441234 706758 441854 711590
rect 441234 706202 441266 706758
rect 441822 706202 441854 706758
rect 441234 694894 441854 706202
rect 441234 694338 441266 694894
rect 441822 694338 441854 694894
rect 441234 658894 441854 694338
rect 441234 658338 441266 658894
rect 441822 658338 441854 658894
rect 441234 622894 441854 658338
rect 441234 622338 441266 622894
rect 441822 622338 441854 622894
rect 441234 586894 441854 622338
rect 441234 586338 441266 586894
rect 441822 586338 441854 586894
rect 441234 550894 441854 586338
rect 441234 550338 441266 550894
rect 441822 550338 441854 550894
rect 441234 514894 441854 550338
rect 441234 514338 441266 514894
rect 441822 514338 441854 514894
rect 441234 478894 441854 514338
rect 441234 478338 441266 478894
rect 441822 478338 441854 478894
rect 441234 442894 441854 478338
rect 441234 442338 441266 442894
rect 441822 442338 441854 442894
rect 441234 406894 441854 442338
rect 441234 406338 441266 406894
rect 441822 406338 441854 406894
rect 441234 370894 441854 406338
rect 441234 370338 441266 370894
rect 441822 370338 441854 370894
rect 441234 334894 441854 370338
rect 441234 334338 441266 334894
rect 441822 334338 441854 334894
rect 441234 298894 441854 334338
rect 441234 298338 441266 298894
rect 441822 298338 441854 298894
rect 441234 262894 441854 298338
rect 441234 262338 441266 262894
rect 441822 262338 441854 262894
rect 441234 226894 441854 262338
rect 441234 226338 441266 226894
rect 441822 226338 441854 226894
rect 441234 190894 441854 226338
rect 441234 190338 441266 190894
rect 441822 190338 441854 190894
rect 441234 154894 441854 190338
rect 441234 154338 441266 154894
rect 441822 154338 441854 154894
rect 441234 118894 441854 154338
rect 441234 118338 441266 118894
rect 441822 118338 441854 118894
rect 441234 82894 441854 118338
rect 441234 82338 441266 82894
rect 441822 82338 441854 82894
rect 441234 46894 441854 82338
rect 441234 46338 441266 46894
rect 441822 46338 441854 46894
rect 441234 10894 441854 46338
rect 441234 10338 441266 10894
rect 441822 10338 441854 10894
rect 441234 -2266 441854 10338
rect 441234 -2822 441266 -2266
rect 441822 -2822 441854 -2266
rect 441234 -7654 441854 -2822
rect 444954 707718 445574 711590
rect 444954 707162 444986 707718
rect 445542 707162 445574 707718
rect 444954 698614 445574 707162
rect 444954 698058 444986 698614
rect 445542 698058 445574 698614
rect 444954 662614 445574 698058
rect 444954 662058 444986 662614
rect 445542 662058 445574 662614
rect 444954 626614 445574 662058
rect 444954 626058 444986 626614
rect 445542 626058 445574 626614
rect 444954 590614 445574 626058
rect 444954 590058 444986 590614
rect 445542 590058 445574 590614
rect 444954 554614 445574 590058
rect 444954 554058 444986 554614
rect 445542 554058 445574 554614
rect 444954 518614 445574 554058
rect 444954 518058 444986 518614
rect 445542 518058 445574 518614
rect 444954 482614 445574 518058
rect 444954 482058 444986 482614
rect 445542 482058 445574 482614
rect 444954 446614 445574 482058
rect 444954 446058 444986 446614
rect 445542 446058 445574 446614
rect 444954 410614 445574 446058
rect 444954 410058 444986 410614
rect 445542 410058 445574 410614
rect 444954 374614 445574 410058
rect 444954 374058 444986 374614
rect 445542 374058 445574 374614
rect 444954 338614 445574 374058
rect 444954 338058 444986 338614
rect 445542 338058 445574 338614
rect 444954 302614 445574 338058
rect 444954 302058 444986 302614
rect 445542 302058 445574 302614
rect 444954 266614 445574 302058
rect 444954 266058 444986 266614
rect 445542 266058 445574 266614
rect 444954 230614 445574 266058
rect 444954 230058 444986 230614
rect 445542 230058 445574 230614
rect 444954 194614 445574 230058
rect 444954 194058 444986 194614
rect 445542 194058 445574 194614
rect 444954 158614 445574 194058
rect 444954 158058 444986 158614
rect 445542 158058 445574 158614
rect 444954 122614 445574 158058
rect 444954 122058 444986 122614
rect 445542 122058 445574 122614
rect 444954 86614 445574 122058
rect 444954 86058 444986 86614
rect 445542 86058 445574 86614
rect 444954 50614 445574 86058
rect 444954 50058 444986 50614
rect 445542 50058 445574 50614
rect 444954 14614 445574 50058
rect 444954 14058 444986 14614
rect 445542 14058 445574 14614
rect 444954 -3226 445574 14058
rect 444954 -3782 444986 -3226
rect 445542 -3782 445574 -3226
rect 444954 -7654 445574 -3782
rect 448674 708678 449294 711590
rect 448674 708122 448706 708678
rect 449262 708122 449294 708678
rect 448674 666334 449294 708122
rect 448674 665778 448706 666334
rect 449262 665778 449294 666334
rect 448674 630334 449294 665778
rect 448674 629778 448706 630334
rect 449262 629778 449294 630334
rect 448674 594334 449294 629778
rect 448674 593778 448706 594334
rect 449262 593778 449294 594334
rect 448674 558334 449294 593778
rect 448674 557778 448706 558334
rect 449262 557778 449294 558334
rect 448674 522334 449294 557778
rect 448674 521778 448706 522334
rect 449262 521778 449294 522334
rect 448674 486334 449294 521778
rect 448674 485778 448706 486334
rect 449262 485778 449294 486334
rect 448674 450334 449294 485778
rect 448674 449778 448706 450334
rect 449262 449778 449294 450334
rect 448674 414334 449294 449778
rect 448674 413778 448706 414334
rect 449262 413778 449294 414334
rect 448674 378334 449294 413778
rect 448674 377778 448706 378334
rect 449262 377778 449294 378334
rect 448674 342334 449294 377778
rect 448674 341778 448706 342334
rect 449262 341778 449294 342334
rect 448674 306334 449294 341778
rect 448674 305778 448706 306334
rect 449262 305778 449294 306334
rect 448674 270334 449294 305778
rect 448674 269778 448706 270334
rect 449262 269778 449294 270334
rect 448674 234334 449294 269778
rect 448674 233778 448706 234334
rect 449262 233778 449294 234334
rect 448674 198334 449294 233778
rect 448674 197778 448706 198334
rect 449262 197778 449294 198334
rect 448674 162334 449294 197778
rect 448674 161778 448706 162334
rect 449262 161778 449294 162334
rect 448674 126334 449294 161778
rect 448674 125778 448706 126334
rect 449262 125778 449294 126334
rect 448674 90334 449294 125778
rect 448674 89778 448706 90334
rect 449262 89778 449294 90334
rect 448674 54334 449294 89778
rect 448674 53778 448706 54334
rect 449262 53778 449294 54334
rect 448674 18334 449294 53778
rect 448674 17778 448706 18334
rect 449262 17778 449294 18334
rect 448674 -4186 449294 17778
rect 448674 -4742 448706 -4186
rect 449262 -4742 449294 -4186
rect 448674 -7654 449294 -4742
rect 452394 709638 453014 711590
rect 452394 709082 452426 709638
rect 452982 709082 453014 709638
rect 452394 670054 453014 709082
rect 452394 669498 452426 670054
rect 452982 669498 453014 670054
rect 452394 634054 453014 669498
rect 452394 633498 452426 634054
rect 452982 633498 453014 634054
rect 452394 598054 453014 633498
rect 452394 597498 452426 598054
rect 452982 597498 453014 598054
rect 452394 562054 453014 597498
rect 452394 561498 452426 562054
rect 452982 561498 453014 562054
rect 452394 526054 453014 561498
rect 452394 525498 452426 526054
rect 452982 525498 453014 526054
rect 452394 490054 453014 525498
rect 452394 489498 452426 490054
rect 452982 489498 453014 490054
rect 452394 454054 453014 489498
rect 452394 453498 452426 454054
rect 452982 453498 453014 454054
rect 452394 418054 453014 453498
rect 452394 417498 452426 418054
rect 452982 417498 453014 418054
rect 452394 382054 453014 417498
rect 452394 381498 452426 382054
rect 452982 381498 453014 382054
rect 452394 346054 453014 381498
rect 452394 345498 452426 346054
rect 452982 345498 453014 346054
rect 452394 310054 453014 345498
rect 452394 309498 452426 310054
rect 452982 309498 453014 310054
rect 452394 274054 453014 309498
rect 452394 273498 452426 274054
rect 452982 273498 453014 274054
rect 452394 238054 453014 273498
rect 452394 237498 452426 238054
rect 452982 237498 453014 238054
rect 452394 202054 453014 237498
rect 452394 201498 452426 202054
rect 452982 201498 453014 202054
rect 452394 166054 453014 201498
rect 452394 165498 452426 166054
rect 452982 165498 453014 166054
rect 452394 130054 453014 165498
rect 452394 129498 452426 130054
rect 452982 129498 453014 130054
rect 452394 94054 453014 129498
rect 452394 93498 452426 94054
rect 452982 93498 453014 94054
rect 452394 58054 453014 93498
rect 452394 57498 452426 58054
rect 452982 57498 453014 58054
rect 452394 22054 453014 57498
rect 452394 21498 452426 22054
rect 452982 21498 453014 22054
rect 452394 -5146 453014 21498
rect 452394 -5702 452426 -5146
rect 452982 -5702 453014 -5146
rect 452394 -7654 453014 -5702
rect 456114 710598 456734 711590
rect 456114 710042 456146 710598
rect 456702 710042 456734 710598
rect 456114 673774 456734 710042
rect 456114 673218 456146 673774
rect 456702 673218 456734 673774
rect 456114 637774 456734 673218
rect 456114 637218 456146 637774
rect 456702 637218 456734 637774
rect 456114 601774 456734 637218
rect 456114 601218 456146 601774
rect 456702 601218 456734 601774
rect 456114 565774 456734 601218
rect 456114 565218 456146 565774
rect 456702 565218 456734 565774
rect 456114 529774 456734 565218
rect 456114 529218 456146 529774
rect 456702 529218 456734 529774
rect 456114 493774 456734 529218
rect 456114 493218 456146 493774
rect 456702 493218 456734 493774
rect 456114 457774 456734 493218
rect 456114 457218 456146 457774
rect 456702 457218 456734 457774
rect 456114 421774 456734 457218
rect 456114 421218 456146 421774
rect 456702 421218 456734 421774
rect 456114 385774 456734 421218
rect 456114 385218 456146 385774
rect 456702 385218 456734 385774
rect 456114 349774 456734 385218
rect 456114 349218 456146 349774
rect 456702 349218 456734 349774
rect 456114 313774 456734 349218
rect 456114 313218 456146 313774
rect 456702 313218 456734 313774
rect 456114 277774 456734 313218
rect 456114 277218 456146 277774
rect 456702 277218 456734 277774
rect 456114 241774 456734 277218
rect 456114 241218 456146 241774
rect 456702 241218 456734 241774
rect 456114 205774 456734 241218
rect 456114 205218 456146 205774
rect 456702 205218 456734 205774
rect 456114 169774 456734 205218
rect 456114 169218 456146 169774
rect 456702 169218 456734 169774
rect 456114 133774 456734 169218
rect 456114 133218 456146 133774
rect 456702 133218 456734 133774
rect 456114 97774 456734 133218
rect 456114 97218 456146 97774
rect 456702 97218 456734 97774
rect 456114 61774 456734 97218
rect 456114 61218 456146 61774
rect 456702 61218 456734 61774
rect 456114 25774 456734 61218
rect 456114 25218 456146 25774
rect 456702 25218 456734 25774
rect 456114 -6106 456734 25218
rect 456114 -6662 456146 -6106
rect 456702 -6662 456734 -6106
rect 456114 -7654 456734 -6662
rect 459834 711558 460454 711590
rect 459834 711002 459866 711558
rect 460422 711002 460454 711558
rect 459834 677494 460454 711002
rect 459834 676938 459866 677494
rect 460422 676938 460454 677494
rect 459834 641494 460454 676938
rect 459834 640938 459866 641494
rect 460422 640938 460454 641494
rect 459834 605494 460454 640938
rect 459834 604938 459866 605494
rect 460422 604938 460454 605494
rect 459834 569494 460454 604938
rect 459834 568938 459866 569494
rect 460422 568938 460454 569494
rect 459834 533494 460454 568938
rect 459834 532938 459866 533494
rect 460422 532938 460454 533494
rect 459834 497494 460454 532938
rect 459834 496938 459866 497494
rect 460422 496938 460454 497494
rect 459834 461494 460454 496938
rect 459834 460938 459866 461494
rect 460422 460938 460454 461494
rect 459834 425494 460454 460938
rect 459834 424938 459866 425494
rect 460422 424938 460454 425494
rect 459834 389494 460454 424938
rect 459834 388938 459866 389494
rect 460422 388938 460454 389494
rect 459834 353494 460454 388938
rect 459834 352938 459866 353494
rect 460422 352938 460454 353494
rect 459834 317494 460454 352938
rect 459834 316938 459866 317494
rect 460422 316938 460454 317494
rect 459834 281494 460454 316938
rect 459834 280938 459866 281494
rect 460422 280938 460454 281494
rect 459834 245494 460454 280938
rect 459834 244938 459866 245494
rect 460422 244938 460454 245494
rect 459834 209494 460454 244938
rect 459834 208938 459866 209494
rect 460422 208938 460454 209494
rect 459834 173494 460454 208938
rect 459834 172938 459866 173494
rect 460422 172938 460454 173494
rect 459834 137494 460454 172938
rect 459834 136938 459866 137494
rect 460422 136938 460454 137494
rect 459834 101494 460454 136938
rect 459834 100938 459866 101494
rect 460422 100938 460454 101494
rect 459834 65494 460454 100938
rect 459834 64938 459866 65494
rect 460422 64938 460454 65494
rect 459834 29494 460454 64938
rect 459834 28938 459866 29494
rect 460422 28938 460454 29494
rect 459834 -7066 460454 28938
rect 459834 -7622 459866 -7066
rect 460422 -7622 460454 -7066
rect 459834 -7654 460454 -7622
rect 469794 704838 470414 711590
rect 469794 704282 469826 704838
rect 470382 704282 470414 704838
rect 469794 687454 470414 704282
rect 469794 686898 469826 687454
rect 470382 686898 470414 687454
rect 469794 651454 470414 686898
rect 469794 650898 469826 651454
rect 470382 650898 470414 651454
rect 469794 615454 470414 650898
rect 469794 614898 469826 615454
rect 470382 614898 470414 615454
rect 469794 579454 470414 614898
rect 469794 578898 469826 579454
rect 470382 578898 470414 579454
rect 469794 543454 470414 578898
rect 469794 542898 469826 543454
rect 470382 542898 470414 543454
rect 469794 507454 470414 542898
rect 469794 506898 469826 507454
rect 470382 506898 470414 507454
rect 469794 471454 470414 506898
rect 469794 470898 469826 471454
rect 470382 470898 470414 471454
rect 469794 435454 470414 470898
rect 469794 434898 469826 435454
rect 470382 434898 470414 435454
rect 469794 399454 470414 434898
rect 469794 398898 469826 399454
rect 470382 398898 470414 399454
rect 469794 363454 470414 398898
rect 469794 362898 469826 363454
rect 470382 362898 470414 363454
rect 469794 327454 470414 362898
rect 469794 326898 469826 327454
rect 470382 326898 470414 327454
rect 469794 291454 470414 326898
rect 469794 290898 469826 291454
rect 470382 290898 470414 291454
rect 469794 255454 470414 290898
rect 469794 254898 469826 255454
rect 470382 254898 470414 255454
rect 469794 219454 470414 254898
rect 469794 218898 469826 219454
rect 470382 218898 470414 219454
rect 469794 183454 470414 218898
rect 469794 182898 469826 183454
rect 470382 182898 470414 183454
rect 469794 147454 470414 182898
rect 469794 146898 469826 147454
rect 470382 146898 470414 147454
rect 469794 111454 470414 146898
rect 469794 110898 469826 111454
rect 470382 110898 470414 111454
rect 469794 75454 470414 110898
rect 469794 74898 469826 75454
rect 470382 74898 470414 75454
rect 469794 39454 470414 74898
rect 469794 38898 469826 39454
rect 470382 38898 470414 39454
rect 469794 3454 470414 38898
rect 469794 2898 469826 3454
rect 470382 2898 470414 3454
rect 469794 -346 470414 2898
rect 469794 -902 469826 -346
rect 470382 -902 470414 -346
rect 469794 -7654 470414 -902
rect 473514 705798 474134 711590
rect 473514 705242 473546 705798
rect 474102 705242 474134 705798
rect 473514 691174 474134 705242
rect 473514 690618 473546 691174
rect 474102 690618 474134 691174
rect 473514 655174 474134 690618
rect 473514 654618 473546 655174
rect 474102 654618 474134 655174
rect 473514 619174 474134 654618
rect 473514 618618 473546 619174
rect 474102 618618 474134 619174
rect 473514 583174 474134 618618
rect 473514 582618 473546 583174
rect 474102 582618 474134 583174
rect 473514 547174 474134 582618
rect 473514 546618 473546 547174
rect 474102 546618 474134 547174
rect 473514 511174 474134 546618
rect 473514 510618 473546 511174
rect 474102 510618 474134 511174
rect 473514 475174 474134 510618
rect 473514 474618 473546 475174
rect 474102 474618 474134 475174
rect 473514 439174 474134 474618
rect 473514 438618 473546 439174
rect 474102 438618 474134 439174
rect 473514 403174 474134 438618
rect 473514 402618 473546 403174
rect 474102 402618 474134 403174
rect 473514 367174 474134 402618
rect 473514 366618 473546 367174
rect 474102 366618 474134 367174
rect 473514 331174 474134 366618
rect 473514 330618 473546 331174
rect 474102 330618 474134 331174
rect 473514 295174 474134 330618
rect 473514 294618 473546 295174
rect 474102 294618 474134 295174
rect 473514 259174 474134 294618
rect 473514 258618 473546 259174
rect 474102 258618 474134 259174
rect 473514 223174 474134 258618
rect 473514 222618 473546 223174
rect 474102 222618 474134 223174
rect 473514 187174 474134 222618
rect 473514 186618 473546 187174
rect 474102 186618 474134 187174
rect 473514 151174 474134 186618
rect 473514 150618 473546 151174
rect 474102 150618 474134 151174
rect 473514 115174 474134 150618
rect 473514 114618 473546 115174
rect 474102 114618 474134 115174
rect 473514 79174 474134 114618
rect 473514 78618 473546 79174
rect 474102 78618 474134 79174
rect 473514 43174 474134 78618
rect 473514 42618 473546 43174
rect 474102 42618 474134 43174
rect 473514 7174 474134 42618
rect 473514 6618 473546 7174
rect 474102 6618 474134 7174
rect 473514 -1306 474134 6618
rect 473514 -1862 473546 -1306
rect 474102 -1862 474134 -1306
rect 473514 -7654 474134 -1862
rect 477234 706758 477854 711590
rect 477234 706202 477266 706758
rect 477822 706202 477854 706758
rect 477234 694894 477854 706202
rect 477234 694338 477266 694894
rect 477822 694338 477854 694894
rect 477234 658894 477854 694338
rect 477234 658338 477266 658894
rect 477822 658338 477854 658894
rect 477234 622894 477854 658338
rect 477234 622338 477266 622894
rect 477822 622338 477854 622894
rect 477234 586894 477854 622338
rect 477234 586338 477266 586894
rect 477822 586338 477854 586894
rect 477234 550894 477854 586338
rect 477234 550338 477266 550894
rect 477822 550338 477854 550894
rect 477234 514894 477854 550338
rect 477234 514338 477266 514894
rect 477822 514338 477854 514894
rect 477234 478894 477854 514338
rect 477234 478338 477266 478894
rect 477822 478338 477854 478894
rect 477234 442894 477854 478338
rect 477234 442338 477266 442894
rect 477822 442338 477854 442894
rect 477234 406894 477854 442338
rect 477234 406338 477266 406894
rect 477822 406338 477854 406894
rect 477234 370894 477854 406338
rect 477234 370338 477266 370894
rect 477822 370338 477854 370894
rect 477234 334894 477854 370338
rect 477234 334338 477266 334894
rect 477822 334338 477854 334894
rect 477234 298894 477854 334338
rect 477234 298338 477266 298894
rect 477822 298338 477854 298894
rect 477234 262894 477854 298338
rect 477234 262338 477266 262894
rect 477822 262338 477854 262894
rect 477234 226894 477854 262338
rect 477234 226338 477266 226894
rect 477822 226338 477854 226894
rect 477234 190894 477854 226338
rect 477234 190338 477266 190894
rect 477822 190338 477854 190894
rect 477234 154894 477854 190338
rect 477234 154338 477266 154894
rect 477822 154338 477854 154894
rect 477234 118894 477854 154338
rect 477234 118338 477266 118894
rect 477822 118338 477854 118894
rect 477234 82894 477854 118338
rect 477234 82338 477266 82894
rect 477822 82338 477854 82894
rect 477234 46894 477854 82338
rect 477234 46338 477266 46894
rect 477822 46338 477854 46894
rect 477234 10894 477854 46338
rect 477234 10338 477266 10894
rect 477822 10338 477854 10894
rect 477234 -2266 477854 10338
rect 477234 -2822 477266 -2266
rect 477822 -2822 477854 -2266
rect 477234 -7654 477854 -2822
rect 480954 707718 481574 711590
rect 480954 707162 480986 707718
rect 481542 707162 481574 707718
rect 480954 698614 481574 707162
rect 480954 698058 480986 698614
rect 481542 698058 481574 698614
rect 480954 662614 481574 698058
rect 480954 662058 480986 662614
rect 481542 662058 481574 662614
rect 480954 626614 481574 662058
rect 480954 626058 480986 626614
rect 481542 626058 481574 626614
rect 480954 590614 481574 626058
rect 480954 590058 480986 590614
rect 481542 590058 481574 590614
rect 480954 554614 481574 590058
rect 480954 554058 480986 554614
rect 481542 554058 481574 554614
rect 480954 518614 481574 554058
rect 480954 518058 480986 518614
rect 481542 518058 481574 518614
rect 480954 482614 481574 518058
rect 480954 482058 480986 482614
rect 481542 482058 481574 482614
rect 480954 446614 481574 482058
rect 480954 446058 480986 446614
rect 481542 446058 481574 446614
rect 480954 410614 481574 446058
rect 480954 410058 480986 410614
rect 481542 410058 481574 410614
rect 480954 374614 481574 410058
rect 480954 374058 480986 374614
rect 481542 374058 481574 374614
rect 480954 338614 481574 374058
rect 480954 338058 480986 338614
rect 481542 338058 481574 338614
rect 480954 302614 481574 338058
rect 480954 302058 480986 302614
rect 481542 302058 481574 302614
rect 480954 266614 481574 302058
rect 480954 266058 480986 266614
rect 481542 266058 481574 266614
rect 480954 230614 481574 266058
rect 480954 230058 480986 230614
rect 481542 230058 481574 230614
rect 480954 194614 481574 230058
rect 480954 194058 480986 194614
rect 481542 194058 481574 194614
rect 480954 158614 481574 194058
rect 480954 158058 480986 158614
rect 481542 158058 481574 158614
rect 480954 122614 481574 158058
rect 480954 122058 480986 122614
rect 481542 122058 481574 122614
rect 480954 86614 481574 122058
rect 480954 86058 480986 86614
rect 481542 86058 481574 86614
rect 480954 50614 481574 86058
rect 480954 50058 480986 50614
rect 481542 50058 481574 50614
rect 480954 14614 481574 50058
rect 480954 14058 480986 14614
rect 481542 14058 481574 14614
rect 480954 -3226 481574 14058
rect 480954 -3782 480986 -3226
rect 481542 -3782 481574 -3226
rect 480954 -7654 481574 -3782
rect 484674 708678 485294 711590
rect 484674 708122 484706 708678
rect 485262 708122 485294 708678
rect 484674 666334 485294 708122
rect 484674 665778 484706 666334
rect 485262 665778 485294 666334
rect 484674 630334 485294 665778
rect 484674 629778 484706 630334
rect 485262 629778 485294 630334
rect 484674 594334 485294 629778
rect 484674 593778 484706 594334
rect 485262 593778 485294 594334
rect 484674 558334 485294 593778
rect 484674 557778 484706 558334
rect 485262 557778 485294 558334
rect 484674 522334 485294 557778
rect 484674 521778 484706 522334
rect 485262 521778 485294 522334
rect 484674 486334 485294 521778
rect 484674 485778 484706 486334
rect 485262 485778 485294 486334
rect 484674 450334 485294 485778
rect 484674 449778 484706 450334
rect 485262 449778 485294 450334
rect 484674 414334 485294 449778
rect 484674 413778 484706 414334
rect 485262 413778 485294 414334
rect 484674 378334 485294 413778
rect 484674 377778 484706 378334
rect 485262 377778 485294 378334
rect 484674 342334 485294 377778
rect 484674 341778 484706 342334
rect 485262 341778 485294 342334
rect 484674 306334 485294 341778
rect 484674 305778 484706 306334
rect 485262 305778 485294 306334
rect 484674 270334 485294 305778
rect 484674 269778 484706 270334
rect 485262 269778 485294 270334
rect 484674 234334 485294 269778
rect 484674 233778 484706 234334
rect 485262 233778 485294 234334
rect 484674 198334 485294 233778
rect 484674 197778 484706 198334
rect 485262 197778 485294 198334
rect 484674 162334 485294 197778
rect 484674 161778 484706 162334
rect 485262 161778 485294 162334
rect 484674 126334 485294 161778
rect 484674 125778 484706 126334
rect 485262 125778 485294 126334
rect 484674 90334 485294 125778
rect 484674 89778 484706 90334
rect 485262 89778 485294 90334
rect 484674 54334 485294 89778
rect 484674 53778 484706 54334
rect 485262 53778 485294 54334
rect 484674 18334 485294 53778
rect 484674 17778 484706 18334
rect 485262 17778 485294 18334
rect 484674 -4186 485294 17778
rect 484674 -4742 484706 -4186
rect 485262 -4742 485294 -4186
rect 484674 -7654 485294 -4742
rect 488394 709638 489014 711590
rect 488394 709082 488426 709638
rect 488982 709082 489014 709638
rect 488394 670054 489014 709082
rect 488394 669498 488426 670054
rect 488982 669498 489014 670054
rect 488394 634054 489014 669498
rect 488394 633498 488426 634054
rect 488982 633498 489014 634054
rect 488394 598054 489014 633498
rect 488394 597498 488426 598054
rect 488982 597498 489014 598054
rect 488394 562054 489014 597498
rect 488394 561498 488426 562054
rect 488982 561498 489014 562054
rect 488394 526054 489014 561498
rect 488394 525498 488426 526054
rect 488982 525498 489014 526054
rect 488394 490054 489014 525498
rect 488394 489498 488426 490054
rect 488982 489498 489014 490054
rect 488394 454054 489014 489498
rect 488394 453498 488426 454054
rect 488982 453498 489014 454054
rect 488394 418054 489014 453498
rect 488394 417498 488426 418054
rect 488982 417498 489014 418054
rect 488394 382054 489014 417498
rect 488394 381498 488426 382054
rect 488982 381498 489014 382054
rect 488394 346054 489014 381498
rect 488394 345498 488426 346054
rect 488982 345498 489014 346054
rect 488394 310054 489014 345498
rect 488394 309498 488426 310054
rect 488982 309498 489014 310054
rect 488394 274054 489014 309498
rect 488394 273498 488426 274054
rect 488982 273498 489014 274054
rect 488394 238054 489014 273498
rect 488394 237498 488426 238054
rect 488982 237498 489014 238054
rect 488394 202054 489014 237498
rect 488394 201498 488426 202054
rect 488982 201498 489014 202054
rect 488394 166054 489014 201498
rect 488394 165498 488426 166054
rect 488982 165498 489014 166054
rect 488394 130054 489014 165498
rect 488394 129498 488426 130054
rect 488982 129498 489014 130054
rect 488394 94054 489014 129498
rect 488394 93498 488426 94054
rect 488982 93498 489014 94054
rect 488394 58054 489014 93498
rect 488394 57498 488426 58054
rect 488982 57498 489014 58054
rect 488394 22054 489014 57498
rect 488394 21498 488426 22054
rect 488982 21498 489014 22054
rect 488394 -5146 489014 21498
rect 488394 -5702 488426 -5146
rect 488982 -5702 489014 -5146
rect 488394 -7654 489014 -5702
rect 492114 710598 492734 711590
rect 492114 710042 492146 710598
rect 492702 710042 492734 710598
rect 492114 673774 492734 710042
rect 492114 673218 492146 673774
rect 492702 673218 492734 673774
rect 492114 637774 492734 673218
rect 492114 637218 492146 637774
rect 492702 637218 492734 637774
rect 492114 601774 492734 637218
rect 492114 601218 492146 601774
rect 492702 601218 492734 601774
rect 492114 565774 492734 601218
rect 492114 565218 492146 565774
rect 492702 565218 492734 565774
rect 492114 529774 492734 565218
rect 492114 529218 492146 529774
rect 492702 529218 492734 529774
rect 492114 493774 492734 529218
rect 492114 493218 492146 493774
rect 492702 493218 492734 493774
rect 492114 457774 492734 493218
rect 492114 457218 492146 457774
rect 492702 457218 492734 457774
rect 492114 421774 492734 457218
rect 492114 421218 492146 421774
rect 492702 421218 492734 421774
rect 492114 385774 492734 421218
rect 492114 385218 492146 385774
rect 492702 385218 492734 385774
rect 492114 349774 492734 385218
rect 492114 349218 492146 349774
rect 492702 349218 492734 349774
rect 492114 313774 492734 349218
rect 492114 313218 492146 313774
rect 492702 313218 492734 313774
rect 492114 277774 492734 313218
rect 492114 277218 492146 277774
rect 492702 277218 492734 277774
rect 492114 241774 492734 277218
rect 492114 241218 492146 241774
rect 492702 241218 492734 241774
rect 492114 205774 492734 241218
rect 492114 205218 492146 205774
rect 492702 205218 492734 205774
rect 492114 169774 492734 205218
rect 492114 169218 492146 169774
rect 492702 169218 492734 169774
rect 492114 133774 492734 169218
rect 492114 133218 492146 133774
rect 492702 133218 492734 133774
rect 492114 97774 492734 133218
rect 492114 97218 492146 97774
rect 492702 97218 492734 97774
rect 492114 61774 492734 97218
rect 492114 61218 492146 61774
rect 492702 61218 492734 61774
rect 492114 25774 492734 61218
rect 492114 25218 492146 25774
rect 492702 25218 492734 25774
rect 492114 -6106 492734 25218
rect 492114 -6662 492146 -6106
rect 492702 -6662 492734 -6106
rect 492114 -7654 492734 -6662
rect 495834 711558 496454 711590
rect 495834 711002 495866 711558
rect 496422 711002 496454 711558
rect 495834 677494 496454 711002
rect 495834 676938 495866 677494
rect 496422 676938 496454 677494
rect 495834 641494 496454 676938
rect 495834 640938 495866 641494
rect 496422 640938 496454 641494
rect 495834 605494 496454 640938
rect 495834 604938 495866 605494
rect 496422 604938 496454 605494
rect 495834 569494 496454 604938
rect 495834 568938 495866 569494
rect 496422 568938 496454 569494
rect 495834 533494 496454 568938
rect 495834 532938 495866 533494
rect 496422 532938 496454 533494
rect 495834 497494 496454 532938
rect 495834 496938 495866 497494
rect 496422 496938 496454 497494
rect 495834 461494 496454 496938
rect 495834 460938 495866 461494
rect 496422 460938 496454 461494
rect 495834 425494 496454 460938
rect 495834 424938 495866 425494
rect 496422 424938 496454 425494
rect 495834 389494 496454 424938
rect 495834 388938 495866 389494
rect 496422 388938 496454 389494
rect 495834 353494 496454 388938
rect 495834 352938 495866 353494
rect 496422 352938 496454 353494
rect 495834 317494 496454 352938
rect 495834 316938 495866 317494
rect 496422 316938 496454 317494
rect 495834 281494 496454 316938
rect 495834 280938 495866 281494
rect 496422 280938 496454 281494
rect 495834 245494 496454 280938
rect 495834 244938 495866 245494
rect 496422 244938 496454 245494
rect 495834 209494 496454 244938
rect 495834 208938 495866 209494
rect 496422 208938 496454 209494
rect 495834 173494 496454 208938
rect 495834 172938 495866 173494
rect 496422 172938 496454 173494
rect 495834 137494 496454 172938
rect 495834 136938 495866 137494
rect 496422 136938 496454 137494
rect 495834 101494 496454 136938
rect 495834 100938 495866 101494
rect 496422 100938 496454 101494
rect 495834 65494 496454 100938
rect 495834 64938 495866 65494
rect 496422 64938 496454 65494
rect 495834 29494 496454 64938
rect 495834 28938 495866 29494
rect 496422 28938 496454 29494
rect 495834 -7066 496454 28938
rect 495834 -7622 495866 -7066
rect 496422 -7622 496454 -7066
rect 495834 -7654 496454 -7622
rect 505794 704838 506414 711590
rect 505794 704282 505826 704838
rect 506382 704282 506414 704838
rect 505794 687454 506414 704282
rect 505794 686898 505826 687454
rect 506382 686898 506414 687454
rect 505794 651454 506414 686898
rect 505794 650898 505826 651454
rect 506382 650898 506414 651454
rect 505794 615454 506414 650898
rect 505794 614898 505826 615454
rect 506382 614898 506414 615454
rect 505794 579454 506414 614898
rect 505794 578898 505826 579454
rect 506382 578898 506414 579454
rect 505794 543454 506414 578898
rect 505794 542898 505826 543454
rect 506382 542898 506414 543454
rect 505794 507454 506414 542898
rect 505794 506898 505826 507454
rect 506382 506898 506414 507454
rect 505794 471454 506414 506898
rect 505794 470898 505826 471454
rect 506382 470898 506414 471454
rect 505794 435454 506414 470898
rect 505794 434898 505826 435454
rect 506382 434898 506414 435454
rect 505794 399454 506414 434898
rect 505794 398898 505826 399454
rect 506382 398898 506414 399454
rect 505794 363454 506414 398898
rect 505794 362898 505826 363454
rect 506382 362898 506414 363454
rect 505794 327454 506414 362898
rect 505794 326898 505826 327454
rect 506382 326898 506414 327454
rect 505794 291454 506414 326898
rect 505794 290898 505826 291454
rect 506382 290898 506414 291454
rect 505794 255454 506414 290898
rect 505794 254898 505826 255454
rect 506382 254898 506414 255454
rect 505794 219454 506414 254898
rect 505794 218898 505826 219454
rect 506382 218898 506414 219454
rect 505794 183454 506414 218898
rect 505794 182898 505826 183454
rect 506382 182898 506414 183454
rect 505794 147454 506414 182898
rect 505794 146898 505826 147454
rect 506382 146898 506414 147454
rect 505794 111454 506414 146898
rect 505794 110898 505826 111454
rect 506382 110898 506414 111454
rect 505794 75454 506414 110898
rect 505794 74898 505826 75454
rect 506382 74898 506414 75454
rect 505794 39454 506414 74898
rect 505794 38898 505826 39454
rect 506382 38898 506414 39454
rect 505794 3454 506414 38898
rect 505794 2898 505826 3454
rect 506382 2898 506414 3454
rect 505794 -346 506414 2898
rect 505794 -902 505826 -346
rect 506382 -902 506414 -346
rect 505794 -7654 506414 -902
rect 509514 705798 510134 711590
rect 509514 705242 509546 705798
rect 510102 705242 510134 705798
rect 509514 691174 510134 705242
rect 509514 690618 509546 691174
rect 510102 690618 510134 691174
rect 509514 655174 510134 690618
rect 509514 654618 509546 655174
rect 510102 654618 510134 655174
rect 509514 619174 510134 654618
rect 509514 618618 509546 619174
rect 510102 618618 510134 619174
rect 509514 583174 510134 618618
rect 509514 582618 509546 583174
rect 510102 582618 510134 583174
rect 509514 547174 510134 582618
rect 509514 546618 509546 547174
rect 510102 546618 510134 547174
rect 509514 511174 510134 546618
rect 509514 510618 509546 511174
rect 510102 510618 510134 511174
rect 509514 475174 510134 510618
rect 509514 474618 509546 475174
rect 510102 474618 510134 475174
rect 509514 439174 510134 474618
rect 509514 438618 509546 439174
rect 510102 438618 510134 439174
rect 509514 403174 510134 438618
rect 509514 402618 509546 403174
rect 510102 402618 510134 403174
rect 509514 367174 510134 402618
rect 509514 366618 509546 367174
rect 510102 366618 510134 367174
rect 509514 331174 510134 366618
rect 509514 330618 509546 331174
rect 510102 330618 510134 331174
rect 509514 295174 510134 330618
rect 509514 294618 509546 295174
rect 510102 294618 510134 295174
rect 509514 259174 510134 294618
rect 509514 258618 509546 259174
rect 510102 258618 510134 259174
rect 509514 223174 510134 258618
rect 509514 222618 509546 223174
rect 510102 222618 510134 223174
rect 509514 187174 510134 222618
rect 509514 186618 509546 187174
rect 510102 186618 510134 187174
rect 509514 151174 510134 186618
rect 509514 150618 509546 151174
rect 510102 150618 510134 151174
rect 509514 115174 510134 150618
rect 509514 114618 509546 115174
rect 510102 114618 510134 115174
rect 509514 79174 510134 114618
rect 509514 78618 509546 79174
rect 510102 78618 510134 79174
rect 509514 43174 510134 78618
rect 509514 42618 509546 43174
rect 510102 42618 510134 43174
rect 509514 7174 510134 42618
rect 509514 6618 509546 7174
rect 510102 6618 510134 7174
rect 509514 -1306 510134 6618
rect 509514 -1862 509546 -1306
rect 510102 -1862 510134 -1306
rect 509514 -7654 510134 -1862
rect 513234 706758 513854 711590
rect 513234 706202 513266 706758
rect 513822 706202 513854 706758
rect 513234 694894 513854 706202
rect 513234 694338 513266 694894
rect 513822 694338 513854 694894
rect 513234 658894 513854 694338
rect 513234 658338 513266 658894
rect 513822 658338 513854 658894
rect 513234 622894 513854 658338
rect 513234 622338 513266 622894
rect 513822 622338 513854 622894
rect 513234 586894 513854 622338
rect 513234 586338 513266 586894
rect 513822 586338 513854 586894
rect 513234 550894 513854 586338
rect 513234 550338 513266 550894
rect 513822 550338 513854 550894
rect 513234 514894 513854 550338
rect 513234 514338 513266 514894
rect 513822 514338 513854 514894
rect 513234 478894 513854 514338
rect 513234 478338 513266 478894
rect 513822 478338 513854 478894
rect 513234 442894 513854 478338
rect 513234 442338 513266 442894
rect 513822 442338 513854 442894
rect 513234 406894 513854 442338
rect 513234 406338 513266 406894
rect 513822 406338 513854 406894
rect 513234 370894 513854 406338
rect 513234 370338 513266 370894
rect 513822 370338 513854 370894
rect 513234 334894 513854 370338
rect 513234 334338 513266 334894
rect 513822 334338 513854 334894
rect 513234 298894 513854 334338
rect 513234 298338 513266 298894
rect 513822 298338 513854 298894
rect 513234 262894 513854 298338
rect 513234 262338 513266 262894
rect 513822 262338 513854 262894
rect 513234 226894 513854 262338
rect 513234 226338 513266 226894
rect 513822 226338 513854 226894
rect 513234 190894 513854 226338
rect 513234 190338 513266 190894
rect 513822 190338 513854 190894
rect 513234 154894 513854 190338
rect 513234 154338 513266 154894
rect 513822 154338 513854 154894
rect 513234 118894 513854 154338
rect 513234 118338 513266 118894
rect 513822 118338 513854 118894
rect 513234 82894 513854 118338
rect 513234 82338 513266 82894
rect 513822 82338 513854 82894
rect 513234 46894 513854 82338
rect 513234 46338 513266 46894
rect 513822 46338 513854 46894
rect 513234 10894 513854 46338
rect 513234 10338 513266 10894
rect 513822 10338 513854 10894
rect 513234 -2266 513854 10338
rect 513234 -2822 513266 -2266
rect 513822 -2822 513854 -2266
rect 513234 -7654 513854 -2822
rect 516954 707718 517574 711590
rect 516954 707162 516986 707718
rect 517542 707162 517574 707718
rect 516954 698614 517574 707162
rect 516954 698058 516986 698614
rect 517542 698058 517574 698614
rect 516954 662614 517574 698058
rect 516954 662058 516986 662614
rect 517542 662058 517574 662614
rect 516954 626614 517574 662058
rect 516954 626058 516986 626614
rect 517542 626058 517574 626614
rect 516954 590614 517574 626058
rect 516954 590058 516986 590614
rect 517542 590058 517574 590614
rect 516954 554614 517574 590058
rect 516954 554058 516986 554614
rect 517542 554058 517574 554614
rect 516954 518614 517574 554058
rect 516954 518058 516986 518614
rect 517542 518058 517574 518614
rect 516954 482614 517574 518058
rect 516954 482058 516986 482614
rect 517542 482058 517574 482614
rect 516954 446614 517574 482058
rect 516954 446058 516986 446614
rect 517542 446058 517574 446614
rect 516954 410614 517574 446058
rect 516954 410058 516986 410614
rect 517542 410058 517574 410614
rect 516954 374614 517574 410058
rect 516954 374058 516986 374614
rect 517542 374058 517574 374614
rect 516954 338614 517574 374058
rect 516954 338058 516986 338614
rect 517542 338058 517574 338614
rect 516954 302614 517574 338058
rect 516954 302058 516986 302614
rect 517542 302058 517574 302614
rect 516954 266614 517574 302058
rect 516954 266058 516986 266614
rect 517542 266058 517574 266614
rect 516954 230614 517574 266058
rect 516954 230058 516986 230614
rect 517542 230058 517574 230614
rect 516954 194614 517574 230058
rect 516954 194058 516986 194614
rect 517542 194058 517574 194614
rect 516954 158614 517574 194058
rect 516954 158058 516986 158614
rect 517542 158058 517574 158614
rect 516954 122614 517574 158058
rect 516954 122058 516986 122614
rect 517542 122058 517574 122614
rect 516954 86614 517574 122058
rect 516954 86058 516986 86614
rect 517542 86058 517574 86614
rect 516954 50614 517574 86058
rect 516954 50058 516986 50614
rect 517542 50058 517574 50614
rect 516954 14614 517574 50058
rect 516954 14058 516986 14614
rect 517542 14058 517574 14614
rect 516954 -3226 517574 14058
rect 516954 -3782 516986 -3226
rect 517542 -3782 517574 -3226
rect 516954 -7654 517574 -3782
rect 520674 708678 521294 711590
rect 520674 708122 520706 708678
rect 521262 708122 521294 708678
rect 520674 666334 521294 708122
rect 520674 665778 520706 666334
rect 521262 665778 521294 666334
rect 520674 630334 521294 665778
rect 520674 629778 520706 630334
rect 521262 629778 521294 630334
rect 520674 594334 521294 629778
rect 520674 593778 520706 594334
rect 521262 593778 521294 594334
rect 520674 558334 521294 593778
rect 520674 557778 520706 558334
rect 521262 557778 521294 558334
rect 520674 522334 521294 557778
rect 520674 521778 520706 522334
rect 521262 521778 521294 522334
rect 520674 486334 521294 521778
rect 520674 485778 520706 486334
rect 521262 485778 521294 486334
rect 520674 450334 521294 485778
rect 520674 449778 520706 450334
rect 521262 449778 521294 450334
rect 520674 414334 521294 449778
rect 520674 413778 520706 414334
rect 521262 413778 521294 414334
rect 520674 378334 521294 413778
rect 520674 377778 520706 378334
rect 521262 377778 521294 378334
rect 520674 342334 521294 377778
rect 520674 341778 520706 342334
rect 521262 341778 521294 342334
rect 520674 306334 521294 341778
rect 520674 305778 520706 306334
rect 521262 305778 521294 306334
rect 520674 270334 521294 305778
rect 520674 269778 520706 270334
rect 521262 269778 521294 270334
rect 520674 234334 521294 269778
rect 520674 233778 520706 234334
rect 521262 233778 521294 234334
rect 520674 198334 521294 233778
rect 520674 197778 520706 198334
rect 521262 197778 521294 198334
rect 520674 162334 521294 197778
rect 520674 161778 520706 162334
rect 521262 161778 521294 162334
rect 520674 126334 521294 161778
rect 520674 125778 520706 126334
rect 521262 125778 521294 126334
rect 520674 90334 521294 125778
rect 520674 89778 520706 90334
rect 521262 89778 521294 90334
rect 520674 54334 521294 89778
rect 520674 53778 520706 54334
rect 521262 53778 521294 54334
rect 520674 18334 521294 53778
rect 520674 17778 520706 18334
rect 521262 17778 521294 18334
rect 520674 -4186 521294 17778
rect 520674 -4742 520706 -4186
rect 521262 -4742 521294 -4186
rect 520674 -7654 521294 -4742
rect 524394 709638 525014 711590
rect 524394 709082 524426 709638
rect 524982 709082 525014 709638
rect 524394 670054 525014 709082
rect 524394 669498 524426 670054
rect 524982 669498 525014 670054
rect 524394 634054 525014 669498
rect 524394 633498 524426 634054
rect 524982 633498 525014 634054
rect 524394 598054 525014 633498
rect 524394 597498 524426 598054
rect 524982 597498 525014 598054
rect 524394 562054 525014 597498
rect 524394 561498 524426 562054
rect 524982 561498 525014 562054
rect 524394 526054 525014 561498
rect 524394 525498 524426 526054
rect 524982 525498 525014 526054
rect 524394 490054 525014 525498
rect 524394 489498 524426 490054
rect 524982 489498 525014 490054
rect 524394 454054 525014 489498
rect 524394 453498 524426 454054
rect 524982 453498 525014 454054
rect 524394 418054 525014 453498
rect 524394 417498 524426 418054
rect 524982 417498 525014 418054
rect 524394 382054 525014 417498
rect 524394 381498 524426 382054
rect 524982 381498 525014 382054
rect 524394 346054 525014 381498
rect 524394 345498 524426 346054
rect 524982 345498 525014 346054
rect 524394 310054 525014 345498
rect 524394 309498 524426 310054
rect 524982 309498 525014 310054
rect 524394 274054 525014 309498
rect 524394 273498 524426 274054
rect 524982 273498 525014 274054
rect 524394 238054 525014 273498
rect 524394 237498 524426 238054
rect 524982 237498 525014 238054
rect 524394 202054 525014 237498
rect 524394 201498 524426 202054
rect 524982 201498 525014 202054
rect 524394 166054 525014 201498
rect 524394 165498 524426 166054
rect 524982 165498 525014 166054
rect 524394 130054 525014 165498
rect 524394 129498 524426 130054
rect 524982 129498 525014 130054
rect 524394 94054 525014 129498
rect 524394 93498 524426 94054
rect 524982 93498 525014 94054
rect 524394 58054 525014 93498
rect 524394 57498 524426 58054
rect 524982 57498 525014 58054
rect 524394 22054 525014 57498
rect 524394 21498 524426 22054
rect 524982 21498 525014 22054
rect 524394 -5146 525014 21498
rect 524394 -5702 524426 -5146
rect 524982 -5702 525014 -5146
rect 524394 -7654 525014 -5702
rect 528114 710598 528734 711590
rect 528114 710042 528146 710598
rect 528702 710042 528734 710598
rect 528114 673774 528734 710042
rect 528114 673218 528146 673774
rect 528702 673218 528734 673774
rect 528114 637774 528734 673218
rect 528114 637218 528146 637774
rect 528702 637218 528734 637774
rect 528114 601774 528734 637218
rect 528114 601218 528146 601774
rect 528702 601218 528734 601774
rect 528114 565774 528734 601218
rect 528114 565218 528146 565774
rect 528702 565218 528734 565774
rect 528114 529774 528734 565218
rect 528114 529218 528146 529774
rect 528702 529218 528734 529774
rect 528114 493774 528734 529218
rect 528114 493218 528146 493774
rect 528702 493218 528734 493774
rect 528114 457774 528734 493218
rect 528114 457218 528146 457774
rect 528702 457218 528734 457774
rect 528114 421774 528734 457218
rect 528114 421218 528146 421774
rect 528702 421218 528734 421774
rect 528114 385774 528734 421218
rect 528114 385218 528146 385774
rect 528702 385218 528734 385774
rect 528114 349774 528734 385218
rect 528114 349218 528146 349774
rect 528702 349218 528734 349774
rect 528114 313774 528734 349218
rect 528114 313218 528146 313774
rect 528702 313218 528734 313774
rect 528114 277774 528734 313218
rect 528114 277218 528146 277774
rect 528702 277218 528734 277774
rect 528114 241774 528734 277218
rect 528114 241218 528146 241774
rect 528702 241218 528734 241774
rect 528114 205774 528734 241218
rect 528114 205218 528146 205774
rect 528702 205218 528734 205774
rect 528114 169774 528734 205218
rect 528114 169218 528146 169774
rect 528702 169218 528734 169774
rect 528114 133774 528734 169218
rect 528114 133218 528146 133774
rect 528702 133218 528734 133774
rect 528114 97774 528734 133218
rect 528114 97218 528146 97774
rect 528702 97218 528734 97774
rect 528114 61774 528734 97218
rect 528114 61218 528146 61774
rect 528702 61218 528734 61774
rect 528114 25774 528734 61218
rect 528114 25218 528146 25774
rect 528702 25218 528734 25774
rect 528114 -6106 528734 25218
rect 528114 -6662 528146 -6106
rect 528702 -6662 528734 -6106
rect 528114 -7654 528734 -6662
rect 531834 711558 532454 711590
rect 531834 711002 531866 711558
rect 532422 711002 532454 711558
rect 531834 677494 532454 711002
rect 531834 676938 531866 677494
rect 532422 676938 532454 677494
rect 531834 641494 532454 676938
rect 531834 640938 531866 641494
rect 532422 640938 532454 641494
rect 531834 605494 532454 640938
rect 531834 604938 531866 605494
rect 532422 604938 532454 605494
rect 531834 569494 532454 604938
rect 531834 568938 531866 569494
rect 532422 568938 532454 569494
rect 531834 533494 532454 568938
rect 531834 532938 531866 533494
rect 532422 532938 532454 533494
rect 531834 497494 532454 532938
rect 531834 496938 531866 497494
rect 532422 496938 532454 497494
rect 531834 461494 532454 496938
rect 531834 460938 531866 461494
rect 532422 460938 532454 461494
rect 531834 425494 532454 460938
rect 531834 424938 531866 425494
rect 532422 424938 532454 425494
rect 531834 389494 532454 424938
rect 531834 388938 531866 389494
rect 532422 388938 532454 389494
rect 531834 353494 532454 388938
rect 531834 352938 531866 353494
rect 532422 352938 532454 353494
rect 531834 317494 532454 352938
rect 531834 316938 531866 317494
rect 532422 316938 532454 317494
rect 531834 281494 532454 316938
rect 531834 280938 531866 281494
rect 532422 280938 532454 281494
rect 531834 245494 532454 280938
rect 531834 244938 531866 245494
rect 532422 244938 532454 245494
rect 531834 209494 532454 244938
rect 531834 208938 531866 209494
rect 532422 208938 532454 209494
rect 531834 173494 532454 208938
rect 531834 172938 531866 173494
rect 532422 172938 532454 173494
rect 531834 137494 532454 172938
rect 531834 136938 531866 137494
rect 532422 136938 532454 137494
rect 531834 101494 532454 136938
rect 531834 100938 531866 101494
rect 532422 100938 532454 101494
rect 531834 65494 532454 100938
rect 531834 64938 531866 65494
rect 532422 64938 532454 65494
rect 531834 29494 532454 64938
rect 531834 28938 531866 29494
rect 532422 28938 532454 29494
rect 531834 -7066 532454 28938
rect 531834 -7622 531866 -7066
rect 532422 -7622 532454 -7066
rect 531834 -7654 532454 -7622
rect 541794 704838 542414 711590
rect 541794 704282 541826 704838
rect 542382 704282 542414 704838
rect 541794 687454 542414 704282
rect 541794 686898 541826 687454
rect 542382 686898 542414 687454
rect 541794 651454 542414 686898
rect 541794 650898 541826 651454
rect 542382 650898 542414 651454
rect 541794 615454 542414 650898
rect 541794 614898 541826 615454
rect 542382 614898 542414 615454
rect 541794 579454 542414 614898
rect 541794 578898 541826 579454
rect 542382 578898 542414 579454
rect 541794 543454 542414 578898
rect 541794 542898 541826 543454
rect 542382 542898 542414 543454
rect 541794 507454 542414 542898
rect 541794 506898 541826 507454
rect 542382 506898 542414 507454
rect 541794 471454 542414 506898
rect 541794 470898 541826 471454
rect 542382 470898 542414 471454
rect 541794 435454 542414 470898
rect 541794 434898 541826 435454
rect 542382 434898 542414 435454
rect 541794 399454 542414 434898
rect 541794 398898 541826 399454
rect 542382 398898 542414 399454
rect 541794 363454 542414 398898
rect 541794 362898 541826 363454
rect 542382 362898 542414 363454
rect 541794 327454 542414 362898
rect 541794 326898 541826 327454
rect 542382 326898 542414 327454
rect 541794 291454 542414 326898
rect 541794 290898 541826 291454
rect 542382 290898 542414 291454
rect 541794 255454 542414 290898
rect 541794 254898 541826 255454
rect 542382 254898 542414 255454
rect 541794 219454 542414 254898
rect 541794 218898 541826 219454
rect 542382 218898 542414 219454
rect 541794 183454 542414 218898
rect 541794 182898 541826 183454
rect 542382 182898 542414 183454
rect 541794 147454 542414 182898
rect 541794 146898 541826 147454
rect 542382 146898 542414 147454
rect 541794 111454 542414 146898
rect 541794 110898 541826 111454
rect 542382 110898 542414 111454
rect 541794 75454 542414 110898
rect 541794 74898 541826 75454
rect 542382 74898 542414 75454
rect 541794 39454 542414 74898
rect 541794 38898 541826 39454
rect 542382 38898 542414 39454
rect 541794 3454 542414 38898
rect 541794 2898 541826 3454
rect 542382 2898 542414 3454
rect 541794 -346 542414 2898
rect 541794 -902 541826 -346
rect 542382 -902 542414 -346
rect 541794 -7654 542414 -902
rect 545514 705798 546134 711590
rect 545514 705242 545546 705798
rect 546102 705242 546134 705798
rect 545514 691174 546134 705242
rect 545514 690618 545546 691174
rect 546102 690618 546134 691174
rect 545514 655174 546134 690618
rect 545514 654618 545546 655174
rect 546102 654618 546134 655174
rect 545514 619174 546134 654618
rect 545514 618618 545546 619174
rect 546102 618618 546134 619174
rect 545514 583174 546134 618618
rect 545514 582618 545546 583174
rect 546102 582618 546134 583174
rect 545514 547174 546134 582618
rect 545514 546618 545546 547174
rect 546102 546618 546134 547174
rect 545514 511174 546134 546618
rect 545514 510618 545546 511174
rect 546102 510618 546134 511174
rect 545514 475174 546134 510618
rect 545514 474618 545546 475174
rect 546102 474618 546134 475174
rect 545514 439174 546134 474618
rect 545514 438618 545546 439174
rect 546102 438618 546134 439174
rect 545514 403174 546134 438618
rect 545514 402618 545546 403174
rect 546102 402618 546134 403174
rect 545514 367174 546134 402618
rect 545514 366618 545546 367174
rect 546102 366618 546134 367174
rect 545514 331174 546134 366618
rect 545514 330618 545546 331174
rect 546102 330618 546134 331174
rect 545514 295174 546134 330618
rect 545514 294618 545546 295174
rect 546102 294618 546134 295174
rect 545514 259174 546134 294618
rect 545514 258618 545546 259174
rect 546102 258618 546134 259174
rect 545514 223174 546134 258618
rect 545514 222618 545546 223174
rect 546102 222618 546134 223174
rect 545514 187174 546134 222618
rect 545514 186618 545546 187174
rect 546102 186618 546134 187174
rect 545514 151174 546134 186618
rect 545514 150618 545546 151174
rect 546102 150618 546134 151174
rect 545514 115174 546134 150618
rect 545514 114618 545546 115174
rect 546102 114618 546134 115174
rect 545514 79174 546134 114618
rect 545514 78618 545546 79174
rect 546102 78618 546134 79174
rect 545514 43174 546134 78618
rect 545514 42618 545546 43174
rect 546102 42618 546134 43174
rect 545514 7174 546134 42618
rect 545514 6618 545546 7174
rect 546102 6618 546134 7174
rect 545514 -1306 546134 6618
rect 545514 -1862 545546 -1306
rect 546102 -1862 546134 -1306
rect 545514 -7654 546134 -1862
rect 549234 706758 549854 711590
rect 549234 706202 549266 706758
rect 549822 706202 549854 706758
rect 549234 694894 549854 706202
rect 549234 694338 549266 694894
rect 549822 694338 549854 694894
rect 549234 658894 549854 694338
rect 549234 658338 549266 658894
rect 549822 658338 549854 658894
rect 549234 622894 549854 658338
rect 549234 622338 549266 622894
rect 549822 622338 549854 622894
rect 549234 586894 549854 622338
rect 549234 586338 549266 586894
rect 549822 586338 549854 586894
rect 549234 550894 549854 586338
rect 549234 550338 549266 550894
rect 549822 550338 549854 550894
rect 549234 514894 549854 550338
rect 549234 514338 549266 514894
rect 549822 514338 549854 514894
rect 549234 478894 549854 514338
rect 549234 478338 549266 478894
rect 549822 478338 549854 478894
rect 549234 442894 549854 478338
rect 549234 442338 549266 442894
rect 549822 442338 549854 442894
rect 549234 406894 549854 442338
rect 549234 406338 549266 406894
rect 549822 406338 549854 406894
rect 549234 370894 549854 406338
rect 549234 370338 549266 370894
rect 549822 370338 549854 370894
rect 549234 334894 549854 370338
rect 549234 334338 549266 334894
rect 549822 334338 549854 334894
rect 549234 298894 549854 334338
rect 549234 298338 549266 298894
rect 549822 298338 549854 298894
rect 549234 262894 549854 298338
rect 549234 262338 549266 262894
rect 549822 262338 549854 262894
rect 549234 226894 549854 262338
rect 549234 226338 549266 226894
rect 549822 226338 549854 226894
rect 549234 190894 549854 226338
rect 549234 190338 549266 190894
rect 549822 190338 549854 190894
rect 549234 154894 549854 190338
rect 549234 154338 549266 154894
rect 549822 154338 549854 154894
rect 549234 118894 549854 154338
rect 549234 118338 549266 118894
rect 549822 118338 549854 118894
rect 549234 82894 549854 118338
rect 549234 82338 549266 82894
rect 549822 82338 549854 82894
rect 549234 46894 549854 82338
rect 549234 46338 549266 46894
rect 549822 46338 549854 46894
rect 549234 10894 549854 46338
rect 549234 10338 549266 10894
rect 549822 10338 549854 10894
rect 549234 -2266 549854 10338
rect 549234 -2822 549266 -2266
rect 549822 -2822 549854 -2266
rect 549234 -7654 549854 -2822
rect 552954 707718 553574 711590
rect 552954 707162 552986 707718
rect 553542 707162 553574 707718
rect 552954 698614 553574 707162
rect 552954 698058 552986 698614
rect 553542 698058 553574 698614
rect 552954 662614 553574 698058
rect 552954 662058 552986 662614
rect 553542 662058 553574 662614
rect 552954 626614 553574 662058
rect 552954 626058 552986 626614
rect 553542 626058 553574 626614
rect 552954 590614 553574 626058
rect 552954 590058 552986 590614
rect 553542 590058 553574 590614
rect 552954 554614 553574 590058
rect 552954 554058 552986 554614
rect 553542 554058 553574 554614
rect 552954 518614 553574 554058
rect 552954 518058 552986 518614
rect 553542 518058 553574 518614
rect 552954 482614 553574 518058
rect 552954 482058 552986 482614
rect 553542 482058 553574 482614
rect 552954 446614 553574 482058
rect 552954 446058 552986 446614
rect 553542 446058 553574 446614
rect 552954 410614 553574 446058
rect 552954 410058 552986 410614
rect 553542 410058 553574 410614
rect 552954 374614 553574 410058
rect 552954 374058 552986 374614
rect 553542 374058 553574 374614
rect 552954 338614 553574 374058
rect 552954 338058 552986 338614
rect 553542 338058 553574 338614
rect 552954 302614 553574 338058
rect 552954 302058 552986 302614
rect 553542 302058 553574 302614
rect 552954 266614 553574 302058
rect 552954 266058 552986 266614
rect 553542 266058 553574 266614
rect 552954 230614 553574 266058
rect 552954 230058 552986 230614
rect 553542 230058 553574 230614
rect 552954 194614 553574 230058
rect 552954 194058 552986 194614
rect 553542 194058 553574 194614
rect 552954 158614 553574 194058
rect 552954 158058 552986 158614
rect 553542 158058 553574 158614
rect 552954 122614 553574 158058
rect 552954 122058 552986 122614
rect 553542 122058 553574 122614
rect 552954 86614 553574 122058
rect 552954 86058 552986 86614
rect 553542 86058 553574 86614
rect 552954 50614 553574 86058
rect 552954 50058 552986 50614
rect 553542 50058 553574 50614
rect 552954 14614 553574 50058
rect 552954 14058 552986 14614
rect 553542 14058 553574 14614
rect 552954 -3226 553574 14058
rect 552954 -3782 552986 -3226
rect 553542 -3782 553574 -3226
rect 552954 -7654 553574 -3782
rect 556674 708678 557294 711590
rect 556674 708122 556706 708678
rect 557262 708122 557294 708678
rect 556674 666334 557294 708122
rect 556674 665778 556706 666334
rect 557262 665778 557294 666334
rect 556674 630334 557294 665778
rect 556674 629778 556706 630334
rect 557262 629778 557294 630334
rect 556674 594334 557294 629778
rect 556674 593778 556706 594334
rect 557262 593778 557294 594334
rect 556674 558334 557294 593778
rect 556674 557778 556706 558334
rect 557262 557778 557294 558334
rect 556674 522334 557294 557778
rect 556674 521778 556706 522334
rect 557262 521778 557294 522334
rect 556674 486334 557294 521778
rect 556674 485778 556706 486334
rect 557262 485778 557294 486334
rect 556674 450334 557294 485778
rect 556674 449778 556706 450334
rect 557262 449778 557294 450334
rect 556674 414334 557294 449778
rect 556674 413778 556706 414334
rect 557262 413778 557294 414334
rect 556674 378334 557294 413778
rect 556674 377778 556706 378334
rect 557262 377778 557294 378334
rect 556674 342334 557294 377778
rect 556674 341778 556706 342334
rect 557262 341778 557294 342334
rect 556674 306334 557294 341778
rect 556674 305778 556706 306334
rect 557262 305778 557294 306334
rect 556674 270334 557294 305778
rect 556674 269778 556706 270334
rect 557262 269778 557294 270334
rect 556674 234334 557294 269778
rect 556674 233778 556706 234334
rect 557262 233778 557294 234334
rect 556674 198334 557294 233778
rect 556674 197778 556706 198334
rect 557262 197778 557294 198334
rect 556674 162334 557294 197778
rect 556674 161778 556706 162334
rect 557262 161778 557294 162334
rect 556674 126334 557294 161778
rect 556674 125778 556706 126334
rect 557262 125778 557294 126334
rect 556674 90334 557294 125778
rect 556674 89778 556706 90334
rect 557262 89778 557294 90334
rect 556674 54334 557294 89778
rect 556674 53778 556706 54334
rect 557262 53778 557294 54334
rect 556674 18334 557294 53778
rect 556674 17778 556706 18334
rect 557262 17778 557294 18334
rect 556674 -4186 557294 17778
rect 556674 -4742 556706 -4186
rect 557262 -4742 557294 -4186
rect 556674 -7654 557294 -4742
rect 560394 709638 561014 711590
rect 560394 709082 560426 709638
rect 560982 709082 561014 709638
rect 560394 670054 561014 709082
rect 560394 669498 560426 670054
rect 560982 669498 561014 670054
rect 560394 634054 561014 669498
rect 560394 633498 560426 634054
rect 560982 633498 561014 634054
rect 560394 598054 561014 633498
rect 560394 597498 560426 598054
rect 560982 597498 561014 598054
rect 560394 562054 561014 597498
rect 560394 561498 560426 562054
rect 560982 561498 561014 562054
rect 560394 526054 561014 561498
rect 560394 525498 560426 526054
rect 560982 525498 561014 526054
rect 560394 490054 561014 525498
rect 560394 489498 560426 490054
rect 560982 489498 561014 490054
rect 560394 454054 561014 489498
rect 560394 453498 560426 454054
rect 560982 453498 561014 454054
rect 560394 418054 561014 453498
rect 560394 417498 560426 418054
rect 560982 417498 561014 418054
rect 560394 382054 561014 417498
rect 560394 381498 560426 382054
rect 560982 381498 561014 382054
rect 560394 346054 561014 381498
rect 560394 345498 560426 346054
rect 560982 345498 561014 346054
rect 560394 310054 561014 345498
rect 560394 309498 560426 310054
rect 560982 309498 561014 310054
rect 560394 274054 561014 309498
rect 560394 273498 560426 274054
rect 560982 273498 561014 274054
rect 560394 238054 561014 273498
rect 560394 237498 560426 238054
rect 560982 237498 561014 238054
rect 560394 202054 561014 237498
rect 560394 201498 560426 202054
rect 560982 201498 561014 202054
rect 560394 166054 561014 201498
rect 560394 165498 560426 166054
rect 560982 165498 561014 166054
rect 560394 130054 561014 165498
rect 560394 129498 560426 130054
rect 560982 129498 561014 130054
rect 560394 94054 561014 129498
rect 560394 93498 560426 94054
rect 560982 93498 561014 94054
rect 560394 58054 561014 93498
rect 560394 57498 560426 58054
rect 560982 57498 561014 58054
rect 560394 22054 561014 57498
rect 560394 21498 560426 22054
rect 560982 21498 561014 22054
rect 560394 -5146 561014 21498
rect 560394 -5702 560426 -5146
rect 560982 -5702 561014 -5146
rect 560394 -7654 561014 -5702
rect 564114 710598 564734 711590
rect 564114 710042 564146 710598
rect 564702 710042 564734 710598
rect 564114 673774 564734 710042
rect 564114 673218 564146 673774
rect 564702 673218 564734 673774
rect 564114 637774 564734 673218
rect 564114 637218 564146 637774
rect 564702 637218 564734 637774
rect 564114 601774 564734 637218
rect 564114 601218 564146 601774
rect 564702 601218 564734 601774
rect 564114 565774 564734 601218
rect 564114 565218 564146 565774
rect 564702 565218 564734 565774
rect 564114 529774 564734 565218
rect 564114 529218 564146 529774
rect 564702 529218 564734 529774
rect 564114 493774 564734 529218
rect 564114 493218 564146 493774
rect 564702 493218 564734 493774
rect 564114 457774 564734 493218
rect 564114 457218 564146 457774
rect 564702 457218 564734 457774
rect 564114 421774 564734 457218
rect 564114 421218 564146 421774
rect 564702 421218 564734 421774
rect 564114 385774 564734 421218
rect 564114 385218 564146 385774
rect 564702 385218 564734 385774
rect 564114 349774 564734 385218
rect 564114 349218 564146 349774
rect 564702 349218 564734 349774
rect 564114 313774 564734 349218
rect 564114 313218 564146 313774
rect 564702 313218 564734 313774
rect 564114 277774 564734 313218
rect 564114 277218 564146 277774
rect 564702 277218 564734 277774
rect 564114 241774 564734 277218
rect 564114 241218 564146 241774
rect 564702 241218 564734 241774
rect 564114 205774 564734 241218
rect 564114 205218 564146 205774
rect 564702 205218 564734 205774
rect 564114 169774 564734 205218
rect 564114 169218 564146 169774
rect 564702 169218 564734 169774
rect 564114 133774 564734 169218
rect 564114 133218 564146 133774
rect 564702 133218 564734 133774
rect 564114 97774 564734 133218
rect 564114 97218 564146 97774
rect 564702 97218 564734 97774
rect 564114 61774 564734 97218
rect 564114 61218 564146 61774
rect 564702 61218 564734 61774
rect 564114 25774 564734 61218
rect 564114 25218 564146 25774
rect 564702 25218 564734 25774
rect 564114 -6106 564734 25218
rect 564114 -6662 564146 -6106
rect 564702 -6662 564734 -6106
rect 564114 -7654 564734 -6662
rect 567834 711558 568454 711590
rect 567834 711002 567866 711558
rect 568422 711002 568454 711558
rect 567834 677494 568454 711002
rect 567834 676938 567866 677494
rect 568422 676938 568454 677494
rect 567834 641494 568454 676938
rect 567834 640938 567866 641494
rect 568422 640938 568454 641494
rect 567834 605494 568454 640938
rect 567834 604938 567866 605494
rect 568422 604938 568454 605494
rect 567834 569494 568454 604938
rect 567834 568938 567866 569494
rect 568422 568938 568454 569494
rect 567834 533494 568454 568938
rect 567834 532938 567866 533494
rect 568422 532938 568454 533494
rect 567834 497494 568454 532938
rect 567834 496938 567866 497494
rect 568422 496938 568454 497494
rect 567834 461494 568454 496938
rect 567834 460938 567866 461494
rect 568422 460938 568454 461494
rect 567834 425494 568454 460938
rect 567834 424938 567866 425494
rect 568422 424938 568454 425494
rect 567834 389494 568454 424938
rect 567834 388938 567866 389494
rect 568422 388938 568454 389494
rect 567834 353494 568454 388938
rect 567834 352938 567866 353494
rect 568422 352938 568454 353494
rect 567834 317494 568454 352938
rect 567834 316938 567866 317494
rect 568422 316938 568454 317494
rect 567834 281494 568454 316938
rect 567834 280938 567866 281494
rect 568422 280938 568454 281494
rect 567834 245494 568454 280938
rect 567834 244938 567866 245494
rect 568422 244938 568454 245494
rect 567834 209494 568454 244938
rect 567834 208938 567866 209494
rect 568422 208938 568454 209494
rect 567834 173494 568454 208938
rect 567834 172938 567866 173494
rect 568422 172938 568454 173494
rect 567834 137494 568454 172938
rect 567834 136938 567866 137494
rect 568422 136938 568454 137494
rect 567834 101494 568454 136938
rect 567834 100938 567866 101494
rect 568422 100938 568454 101494
rect 567834 65494 568454 100938
rect 567834 64938 567866 65494
rect 568422 64938 568454 65494
rect 567834 29494 568454 64938
rect 567834 28938 567866 29494
rect 568422 28938 568454 29494
rect 567834 -7066 568454 28938
rect 567834 -7622 567866 -7066
rect 568422 -7622 568454 -7066
rect 567834 -7654 568454 -7622
rect 577794 704838 578414 711590
rect 577794 704282 577826 704838
rect 578382 704282 578414 704838
rect 577794 687454 578414 704282
rect 577794 686898 577826 687454
rect 578382 686898 578414 687454
rect 577794 651454 578414 686898
rect 577794 650898 577826 651454
rect 578382 650898 578414 651454
rect 577794 615454 578414 650898
rect 581514 705798 582134 711590
rect 592030 711558 592650 711590
rect 592030 711002 592062 711558
rect 592618 711002 592650 711558
rect 591070 710598 591690 710630
rect 591070 710042 591102 710598
rect 591658 710042 591690 710598
rect 590110 709638 590730 709670
rect 590110 709082 590142 709638
rect 590698 709082 590730 709638
rect 589150 708678 589770 708710
rect 589150 708122 589182 708678
rect 589738 708122 589770 708678
rect 588190 707718 588810 707750
rect 588190 707162 588222 707718
rect 588778 707162 588810 707718
rect 587230 706758 587850 706790
rect 587230 706202 587262 706758
rect 587818 706202 587850 706758
rect 581514 705242 581546 705798
rect 582102 705242 582134 705798
rect 581514 691174 582134 705242
rect 586270 705798 586890 705830
rect 586270 705242 586302 705798
rect 586858 705242 586890 705798
rect 581514 690618 581546 691174
rect 582102 690618 582134 691174
rect 581514 655174 582134 690618
rect 581514 654618 581546 655174
rect 582102 654618 582134 655174
rect 581514 619174 582134 654618
rect 581514 618618 581546 619174
rect 582102 618618 582134 619174
rect 580395 617540 580461 617541
rect 580395 617476 580396 617540
rect 580460 617476 580461 617540
rect 580395 617475 580461 617476
rect 577794 614898 577826 615454
rect 578382 614898 578414 615454
rect 577794 579454 578414 614898
rect 577794 578898 577826 579454
rect 578382 578898 578414 579454
rect 577794 543454 578414 578898
rect 577794 542898 577826 543454
rect 578382 542898 578414 543454
rect 577794 507454 578414 542898
rect 577794 506898 577826 507454
rect 578382 506898 578414 507454
rect 577794 471454 578414 506898
rect 577794 470898 577826 471454
rect 578382 470898 578414 471454
rect 577794 435454 578414 470898
rect 577794 434898 577826 435454
rect 578382 434898 578414 435454
rect 577794 399454 578414 434898
rect 577794 398898 577826 399454
rect 578382 398898 578414 399454
rect 577794 363454 578414 398898
rect 577794 362898 577826 363454
rect 578382 362898 578414 363454
rect 577794 327454 578414 362898
rect 577794 326898 577826 327454
rect 578382 326898 578414 327454
rect 577794 291454 578414 326898
rect 577794 290898 577826 291454
rect 578382 290898 578414 291454
rect 577794 255454 578414 290898
rect 577794 254898 577826 255454
rect 578382 254898 578414 255454
rect 577794 219454 578414 254898
rect 577794 218898 577826 219454
rect 578382 218898 578414 219454
rect 577794 183454 578414 218898
rect 577794 182898 577826 183454
rect 578382 182898 578414 183454
rect 577794 147454 578414 182898
rect 577794 146898 577826 147454
rect 578382 146898 578414 147454
rect 577794 111454 578414 146898
rect 577794 110898 577826 111454
rect 578382 110898 578414 111454
rect 577794 75454 578414 110898
rect 577794 74898 577826 75454
rect 578382 74898 578414 75454
rect 577794 39454 578414 74898
rect 577794 38898 577826 39454
rect 578382 38898 578414 39454
rect 577794 3454 578414 38898
rect 577794 2898 577826 3454
rect 578382 2898 578414 3454
rect 577794 -346 578414 2898
rect 580398 1325 580458 617475
rect 581514 583174 582134 618618
rect 581514 582618 581546 583174
rect 582102 582618 582134 583174
rect 580579 564364 580645 564365
rect 580579 564300 580580 564364
rect 580644 564300 580645 564364
rect 580579 564299 580645 564300
rect 580395 1324 580461 1325
rect 580395 1260 580396 1324
rect 580460 1260 580461 1324
rect 580395 1259 580461 1260
rect 580582 917 580642 564299
rect 581514 547174 582134 582618
rect 581514 546618 581546 547174
rect 582102 546618 582134 547174
rect 581514 511174 582134 546618
rect 581514 510618 581546 511174
rect 582102 510618 582134 511174
rect 581514 475174 582134 510618
rect 581514 474618 581546 475174
rect 582102 474618 582134 475174
rect 581514 439174 582134 474618
rect 581514 438618 581546 439174
rect 582102 438618 582134 439174
rect 581514 403174 582134 438618
rect 581514 402618 581546 403174
rect 582102 402618 582134 403174
rect 581514 367174 582134 402618
rect 581514 366618 581546 367174
rect 582102 366618 582134 367174
rect 581514 331174 582134 366618
rect 581514 330618 581546 331174
rect 582102 330618 582134 331174
rect 581514 295174 582134 330618
rect 581514 294618 581546 295174
rect 582102 294618 582134 295174
rect 581514 259174 582134 294618
rect 581514 258618 581546 259174
rect 582102 258618 582134 259174
rect 581514 223174 582134 258618
rect 581514 222618 581546 223174
rect 582102 222618 582134 223174
rect 581514 187174 582134 222618
rect 581514 186618 581546 187174
rect 582102 186618 582134 187174
rect 581514 151174 582134 186618
rect 581514 150618 581546 151174
rect 582102 150618 582134 151174
rect 581514 115174 582134 150618
rect 581514 114618 581546 115174
rect 582102 114618 582134 115174
rect 581514 79174 582134 114618
rect 581514 78618 581546 79174
rect 582102 78618 582134 79174
rect 581514 43174 582134 78618
rect 581514 42618 581546 43174
rect 582102 42618 582134 43174
rect 581514 7174 582134 42618
rect 581514 6618 581546 7174
rect 582102 6618 582134 7174
rect 580579 916 580645 917
rect 580579 852 580580 916
rect 580644 852 580645 916
rect 580579 851 580645 852
rect 577794 -902 577826 -346
rect 578382 -902 578414 -346
rect 577794 -7654 578414 -902
rect 581514 -1306 582134 6618
rect 585310 704838 585930 704870
rect 585310 704282 585342 704838
rect 585898 704282 585930 704838
rect 585310 687454 585930 704282
rect 585310 686898 585342 687454
rect 585898 686898 585930 687454
rect 585310 651454 585930 686898
rect 585310 650898 585342 651454
rect 585898 650898 585930 651454
rect 585310 615454 585930 650898
rect 585310 614898 585342 615454
rect 585898 614898 585930 615454
rect 585310 579454 585930 614898
rect 585310 578898 585342 579454
rect 585898 578898 585930 579454
rect 585310 543454 585930 578898
rect 585310 542898 585342 543454
rect 585898 542898 585930 543454
rect 585310 507454 585930 542898
rect 585310 506898 585342 507454
rect 585898 506898 585930 507454
rect 585310 471454 585930 506898
rect 585310 470898 585342 471454
rect 585898 470898 585930 471454
rect 585310 435454 585930 470898
rect 585310 434898 585342 435454
rect 585898 434898 585930 435454
rect 585310 399454 585930 434898
rect 585310 398898 585342 399454
rect 585898 398898 585930 399454
rect 585310 363454 585930 398898
rect 585310 362898 585342 363454
rect 585898 362898 585930 363454
rect 585310 327454 585930 362898
rect 585310 326898 585342 327454
rect 585898 326898 585930 327454
rect 585310 291454 585930 326898
rect 585310 290898 585342 291454
rect 585898 290898 585930 291454
rect 585310 255454 585930 290898
rect 585310 254898 585342 255454
rect 585898 254898 585930 255454
rect 585310 219454 585930 254898
rect 585310 218898 585342 219454
rect 585898 218898 585930 219454
rect 585310 183454 585930 218898
rect 585310 182898 585342 183454
rect 585898 182898 585930 183454
rect 585310 147454 585930 182898
rect 585310 146898 585342 147454
rect 585898 146898 585930 147454
rect 585310 111454 585930 146898
rect 585310 110898 585342 111454
rect 585898 110898 585930 111454
rect 585310 75454 585930 110898
rect 585310 74898 585342 75454
rect 585898 74898 585930 75454
rect 585310 39454 585930 74898
rect 585310 38898 585342 39454
rect 585898 38898 585930 39454
rect 585310 3454 585930 38898
rect 585310 2898 585342 3454
rect 585898 2898 585930 3454
rect 585310 -346 585930 2898
rect 585310 -902 585342 -346
rect 585898 -902 585930 -346
rect 585310 -934 585930 -902
rect 586270 691174 586890 705242
rect 586270 690618 586302 691174
rect 586858 690618 586890 691174
rect 586270 655174 586890 690618
rect 586270 654618 586302 655174
rect 586858 654618 586890 655174
rect 586270 619174 586890 654618
rect 586270 618618 586302 619174
rect 586858 618618 586890 619174
rect 586270 583174 586890 618618
rect 586270 582618 586302 583174
rect 586858 582618 586890 583174
rect 586270 547174 586890 582618
rect 586270 546618 586302 547174
rect 586858 546618 586890 547174
rect 586270 511174 586890 546618
rect 586270 510618 586302 511174
rect 586858 510618 586890 511174
rect 586270 475174 586890 510618
rect 586270 474618 586302 475174
rect 586858 474618 586890 475174
rect 586270 439174 586890 474618
rect 586270 438618 586302 439174
rect 586858 438618 586890 439174
rect 586270 403174 586890 438618
rect 586270 402618 586302 403174
rect 586858 402618 586890 403174
rect 586270 367174 586890 402618
rect 586270 366618 586302 367174
rect 586858 366618 586890 367174
rect 586270 331174 586890 366618
rect 586270 330618 586302 331174
rect 586858 330618 586890 331174
rect 586270 295174 586890 330618
rect 586270 294618 586302 295174
rect 586858 294618 586890 295174
rect 586270 259174 586890 294618
rect 586270 258618 586302 259174
rect 586858 258618 586890 259174
rect 586270 223174 586890 258618
rect 586270 222618 586302 223174
rect 586858 222618 586890 223174
rect 586270 187174 586890 222618
rect 586270 186618 586302 187174
rect 586858 186618 586890 187174
rect 586270 151174 586890 186618
rect 586270 150618 586302 151174
rect 586858 150618 586890 151174
rect 586270 115174 586890 150618
rect 586270 114618 586302 115174
rect 586858 114618 586890 115174
rect 586270 79174 586890 114618
rect 586270 78618 586302 79174
rect 586858 78618 586890 79174
rect 586270 43174 586890 78618
rect 586270 42618 586302 43174
rect 586858 42618 586890 43174
rect 586270 7174 586890 42618
rect 586270 6618 586302 7174
rect 586858 6618 586890 7174
rect 581514 -1862 581546 -1306
rect 582102 -1862 582134 -1306
rect 581514 -7654 582134 -1862
rect 586270 -1306 586890 6618
rect 586270 -1862 586302 -1306
rect 586858 -1862 586890 -1306
rect 586270 -1894 586890 -1862
rect 587230 694894 587850 706202
rect 587230 694338 587262 694894
rect 587818 694338 587850 694894
rect 587230 658894 587850 694338
rect 587230 658338 587262 658894
rect 587818 658338 587850 658894
rect 587230 622894 587850 658338
rect 587230 622338 587262 622894
rect 587818 622338 587850 622894
rect 587230 586894 587850 622338
rect 587230 586338 587262 586894
rect 587818 586338 587850 586894
rect 587230 550894 587850 586338
rect 587230 550338 587262 550894
rect 587818 550338 587850 550894
rect 587230 514894 587850 550338
rect 587230 514338 587262 514894
rect 587818 514338 587850 514894
rect 587230 478894 587850 514338
rect 587230 478338 587262 478894
rect 587818 478338 587850 478894
rect 587230 442894 587850 478338
rect 587230 442338 587262 442894
rect 587818 442338 587850 442894
rect 587230 406894 587850 442338
rect 587230 406338 587262 406894
rect 587818 406338 587850 406894
rect 587230 370894 587850 406338
rect 587230 370338 587262 370894
rect 587818 370338 587850 370894
rect 587230 334894 587850 370338
rect 587230 334338 587262 334894
rect 587818 334338 587850 334894
rect 587230 298894 587850 334338
rect 587230 298338 587262 298894
rect 587818 298338 587850 298894
rect 587230 262894 587850 298338
rect 587230 262338 587262 262894
rect 587818 262338 587850 262894
rect 587230 226894 587850 262338
rect 587230 226338 587262 226894
rect 587818 226338 587850 226894
rect 587230 190894 587850 226338
rect 587230 190338 587262 190894
rect 587818 190338 587850 190894
rect 587230 154894 587850 190338
rect 587230 154338 587262 154894
rect 587818 154338 587850 154894
rect 587230 118894 587850 154338
rect 587230 118338 587262 118894
rect 587818 118338 587850 118894
rect 587230 82894 587850 118338
rect 587230 82338 587262 82894
rect 587818 82338 587850 82894
rect 587230 46894 587850 82338
rect 587230 46338 587262 46894
rect 587818 46338 587850 46894
rect 587230 10894 587850 46338
rect 587230 10338 587262 10894
rect 587818 10338 587850 10894
rect 587230 -2266 587850 10338
rect 587230 -2822 587262 -2266
rect 587818 -2822 587850 -2266
rect 587230 -2854 587850 -2822
rect 588190 698614 588810 707162
rect 588190 698058 588222 698614
rect 588778 698058 588810 698614
rect 588190 662614 588810 698058
rect 588190 662058 588222 662614
rect 588778 662058 588810 662614
rect 588190 626614 588810 662058
rect 588190 626058 588222 626614
rect 588778 626058 588810 626614
rect 588190 590614 588810 626058
rect 588190 590058 588222 590614
rect 588778 590058 588810 590614
rect 588190 554614 588810 590058
rect 588190 554058 588222 554614
rect 588778 554058 588810 554614
rect 588190 518614 588810 554058
rect 588190 518058 588222 518614
rect 588778 518058 588810 518614
rect 588190 482614 588810 518058
rect 588190 482058 588222 482614
rect 588778 482058 588810 482614
rect 588190 446614 588810 482058
rect 588190 446058 588222 446614
rect 588778 446058 588810 446614
rect 588190 410614 588810 446058
rect 588190 410058 588222 410614
rect 588778 410058 588810 410614
rect 588190 374614 588810 410058
rect 588190 374058 588222 374614
rect 588778 374058 588810 374614
rect 588190 338614 588810 374058
rect 588190 338058 588222 338614
rect 588778 338058 588810 338614
rect 588190 302614 588810 338058
rect 588190 302058 588222 302614
rect 588778 302058 588810 302614
rect 588190 266614 588810 302058
rect 588190 266058 588222 266614
rect 588778 266058 588810 266614
rect 588190 230614 588810 266058
rect 588190 230058 588222 230614
rect 588778 230058 588810 230614
rect 588190 194614 588810 230058
rect 588190 194058 588222 194614
rect 588778 194058 588810 194614
rect 588190 158614 588810 194058
rect 588190 158058 588222 158614
rect 588778 158058 588810 158614
rect 588190 122614 588810 158058
rect 588190 122058 588222 122614
rect 588778 122058 588810 122614
rect 588190 86614 588810 122058
rect 588190 86058 588222 86614
rect 588778 86058 588810 86614
rect 588190 50614 588810 86058
rect 588190 50058 588222 50614
rect 588778 50058 588810 50614
rect 588190 14614 588810 50058
rect 588190 14058 588222 14614
rect 588778 14058 588810 14614
rect 588190 -3226 588810 14058
rect 588190 -3782 588222 -3226
rect 588778 -3782 588810 -3226
rect 588190 -3814 588810 -3782
rect 589150 666334 589770 708122
rect 589150 665778 589182 666334
rect 589738 665778 589770 666334
rect 589150 630334 589770 665778
rect 589150 629778 589182 630334
rect 589738 629778 589770 630334
rect 589150 594334 589770 629778
rect 589150 593778 589182 594334
rect 589738 593778 589770 594334
rect 589150 558334 589770 593778
rect 589150 557778 589182 558334
rect 589738 557778 589770 558334
rect 589150 522334 589770 557778
rect 589150 521778 589182 522334
rect 589738 521778 589770 522334
rect 589150 486334 589770 521778
rect 589150 485778 589182 486334
rect 589738 485778 589770 486334
rect 589150 450334 589770 485778
rect 589150 449778 589182 450334
rect 589738 449778 589770 450334
rect 589150 414334 589770 449778
rect 589150 413778 589182 414334
rect 589738 413778 589770 414334
rect 589150 378334 589770 413778
rect 589150 377778 589182 378334
rect 589738 377778 589770 378334
rect 589150 342334 589770 377778
rect 589150 341778 589182 342334
rect 589738 341778 589770 342334
rect 589150 306334 589770 341778
rect 589150 305778 589182 306334
rect 589738 305778 589770 306334
rect 589150 270334 589770 305778
rect 589150 269778 589182 270334
rect 589738 269778 589770 270334
rect 589150 234334 589770 269778
rect 589150 233778 589182 234334
rect 589738 233778 589770 234334
rect 589150 198334 589770 233778
rect 589150 197778 589182 198334
rect 589738 197778 589770 198334
rect 589150 162334 589770 197778
rect 589150 161778 589182 162334
rect 589738 161778 589770 162334
rect 589150 126334 589770 161778
rect 589150 125778 589182 126334
rect 589738 125778 589770 126334
rect 589150 90334 589770 125778
rect 589150 89778 589182 90334
rect 589738 89778 589770 90334
rect 589150 54334 589770 89778
rect 589150 53778 589182 54334
rect 589738 53778 589770 54334
rect 589150 18334 589770 53778
rect 589150 17778 589182 18334
rect 589738 17778 589770 18334
rect 589150 -4186 589770 17778
rect 589150 -4742 589182 -4186
rect 589738 -4742 589770 -4186
rect 589150 -4774 589770 -4742
rect 590110 670054 590730 709082
rect 590110 669498 590142 670054
rect 590698 669498 590730 670054
rect 590110 634054 590730 669498
rect 590110 633498 590142 634054
rect 590698 633498 590730 634054
rect 590110 598054 590730 633498
rect 590110 597498 590142 598054
rect 590698 597498 590730 598054
rect 590110 562054 590730 597498
rect 590110 561498 590142 562054
rect 590698 561498 590730 562054
rect 590110 526054 590730 561498
rect 590110 525498 590142 526054
rect 590698 525498 590730 526054
rect 590110 490054 590730 525498
rect 590110 489498 590142 490054
rect 590698 489498 590730 490054
rect 590110 454054 590730 489498
rect 590110 453498 590142 454054
rect 590698 453498 590730 454054
rect 590110 418054 590730 453498
rect 590110 417498 590142 418054
rect 590698 417498 590730 418054
rect 590110 382054 590730 417498
rect 590110 381498 590142 382054
rect 590698 381498 590730 382054
rect 590110 346054 590730 381498
rect 590110 345498 590142 346054
rect 590698 345498 590730 346054
rect 590110 310054 590730 345498
rect 590110 309498 590142 310054
rect 590698 309498 590730 310054
rect 590110 274054 590730 309498
rect 590110 273498 590142 274054
rect 590698 273498 590730 274054
rect 590110 238054 590730 273498
rect 590110 237498 590142 238054
rect 590698 237498 590730 238054
rect 590110 202054 590730 237498
rect 590110 201498 590142 202054
rect 590698 201498 590730 202054
rect 590110 166054 590730 201498
rect 590110 165498 590142 166054
rect 590698 165498 590730 166054
rect 590110 130054 590730 165498
rect 590110 129498 590142 130054
rect 590698 129498 590730 130054
rect 590110 94054 590730 129498
rect 590110 93498 590142 94054
rect 590698 93498 590730 94054
rect 590110 58054 590730 93498
rect 590110 57498 590142 58054
rect 590698 57498 590730 58054
rect 590110 22054 590730 57498
rect 590110 21498 590142 22054
rect 590698 21498 590730 22054
rect 590110 -5146 590730 21498
rect 590110 -5702 590142 -5146
rect 590698 -5702 590730 -5146
rect 590110 -5734 590730 -5702
rect 591070 673774 591690 710042
rect 591070 673218 591102 673774
rect 591658 673218 591690 673774
rect 591070 637774 591690 673218
rect 591070 637218 591102 637774
rect 591658 637218 591690 637774
rect 591070 601774 591690 637218
rect 591070 601218 591102 601774
rect 591658 601218 591690 601774
rect 591070 565774 591690 601218
rect 591070 565218 591102 565774
rect 591658 565218 591690 565774
rect 591070 529774 591690 565218
rect 591070 529218 591102 529774
rect 591658 529218 591690 529774
rect 591070 493774 591690 529218
rect 591070 493218 591102 493774
rect 591658 493218 591690 493774
rect 591070 457774 591690 493218
rect 591070 457218 591102 457774
rect 591658 457218 591690 457774
rect 591070 421774 591690 457218
rect 591070 421218 591102 421774
rect 591658 421218 591690 421774
rect 591070 385774 591690 421218
rect 591070 385218 591102 385774
rect 591658 385218 591690 385774
rect 591070 349774 591690 385218
rect 591070 349218 591102 349774
rect 591658 349218 591690 349774
rect 591070 313774 591690 349218
rect 591070 313218 591102 313774
rect 591658 313218 591690 313774
rect 591070 277774 591690 313218
rect 591070 277218 591102 277774
rect 591658 277218 591690 277774
rect 591070 241774 591690 277218
rect 591070 241218 591102 241774
rect 591658 241218 591690 241774
rect 591070 205774 591690 241218
rect 591070 205218 591102 205774
rect 591658 205218 591690 205774
rect 591070 169774 591690 205218
rect 591070 169218 591102 169774
rect 591658 169218 591690 169774
rect 591070 133774 591690 169218
rect 591070 133218 591102 133774
rect 591658 133218 591690 133774
rect 591070 97774 591690 133218
rect 591070 97218 591102 97774
rect 591658 97218 591690 97774
rect 591070 61774 591690 97218
rect 591070 61218 591102 61774
rect 591658 61218 591690 61774
rect 591070 25774 591690 61218
rect 591070 25218 591102 25774
rect 591658 25218 591690 25774
rect 591070 -6106 591690 25218
rect 591070 -6662 591102 -6106
rect 591658 -6662 591690 -6106
rect 591070 -6694 591690 -6662
rect 592030 677494 592650 711002
rect 592030 676938 592062 677494
rect 592618 676938 592650 677494
rect 592030 641494 592650 676938
rect 592030 640938 592062 641494
rect 592618 640938 592650 641494
rect 592030 605494 592650 640938
rect 592030 604938 592062 605494
rect 592618 604938 592650 605494
rect 592030 569494 592650 604938
rect 592030 568938 592062 569494
rect 592618 568938 592650 569494
rect 592030 533494 592650 568938
rect 592030 532938 592062 533494
rect 592618 532938 592650 533494
rect 592030 497494 592650 532938
rect 592030 496938 592062 497494
rect 592618 496938 592650 497494
rect 592030 461494 592650 496938
rect 592030 460938 592062 461494
rect 592618 460938 592650 461494
rect 592030 425494 592650 460938
rect 592030 424938 592062 425494
rect 592618 424938 592650 425494
rect 592030 389494 592650 424938
rect 592030 388938 592062 389494
rect 592618 388938 592650 389494
rect 592030 353494 592650 388938
rect 592030 352938 592062 353494
rect 592618 352938 592650 353494
rect 592030 317494 592650 352938
rect 592030 316938 592062 317494
rect 592618 316938 592650 317494
rect 592030 281494 592650 316938
rect 592030 280938 592062 281494
rect 592618 280938 592650 281494
rect 592030 245494 592650 280938
rect 592030 244938 592062 245494
rect 592618 244938 592650 245494
rect 592030 209494 592650 244938
rect 592030 208938 592062 209494
rect 592618 208938 592650 209494
rect 592030 173494 592650 208938
rect 592030 172938 592062 173494
rect 592618 172938 592650 173494
rect 592030 137494 592650 172938
rect 592030 136938 592062 137494
rect 592618 136938 592650 137494
rect 592030 101494 592650 136938
rect 592030 100938 592062 101494
rect 592618 100938 592650 101494
rect 592030 65494 592650 100938
rect 592030 64938 592062 65494
rect 592618 64938 592650 65494
rect 592030 29494 592650 64938
rect 592030 28938 592062 29494
rect 592618 28938 592650 29494
rect 592030 -7066 592650 28938
rect 592030 -7622 592062 -7066
rect 592618 -7622 592650 -7066
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711002 -8138 711558
rect -8694 676938 -8138 677494
rect -8694 640938 -8138 641494
rect -8694 604938 -8138 605494
rect -8694 568938 -8138 569494
rect -8694 532938 -8138 533494
rect -8694 496938 -8138 497494
rect -8694 460938 -8138 461494
rect -8694 424938 -8138 425494
rect -8694 388938 -8138 389494
rect -8694 352938 -8138 353494
rect -8694 316938 -8138 317494
rect -8694 280938 -8138 281494
rect -8694 244938 -8138 245494
rect -8694 208938 -8138 209494
rect -8694 172938 -8138 173494
rect -8694 136938 -8138 137494
rect -8694 100938 -8138 101494
rect -8694 64938 -8138 65494
rect -8694 28938 -8138 29494
rect -7734 710042 -7178 710598
rect -7734 673218 -7178 673774
rect -7734 637218 -7178 637774
rect -7734 601218 -7178 601774
rect -7734 565218 -7178 565774
rect -7734 529218 -7178 529774
rect -7734 493218 -7178 493774
rect -7734 457218 -7178 457774
rect -7734 421218 -7178 421774
rect -7734 385218 -7178 385774
rect -7734 349218 -7178 349774
rect -7734 313218 -7178 313774
rect -7734 277218 -7178 277774
rect -7734 241218 -7178 241774
rect -7734 205218 -7178 205774
rect -7734 169218 -7178 169774
rect -7734 133218 -7178 133774
rect -7734 97218 -7178 97774
rect -7734 61218 -7178 61774
rect -7734 25218 -7178 25774
rect -6774 709082 -6218 709638
rect -6774 669498 -6218 670054
rect -6774 633498 -6218 634054
rect -6774 597498 -6218 598054
rect -6774 561498 -6218 562054
rect -6774 525498 -6218 526054
rect -6774 489498 -6218 490054
rect -6774 453498 -6218 454054
rect -6774 417498 -6218 418054
rect -6774 381498 -6218 382054
rect -6774 345498 -6218 346054
rect -6774 309498 -6218 310054
rect -6774 273498 -6218 274054
rect -6774 237498 -6218 238054
rect -6774 201498 -6218 202054
rect -6774 165498 -6218 166054
rect -6774 129498 -6218 130054
rect -6774 93498 -6218 94054
rect -6774 57498 -6218 58054
rect -6774 21498 -6218 22054
rect -5814 708122 -5258 708678
rect -5814 665778 -5258 666334
rect -5814 629778 -5258 630334
rect -5814 593778 -5258 594334
rect -5814 557778 -5258 558334
rect -5814 521778 -5258 522334
rect -5814 485778 -5258 486334
rect -5814 449778 -5258 450334
rect -5814 413778 -5258 414334
rect -5814 377778 -5258 378334
rect -5814 341778 -5258 342334
rect -5814 305778 -5258 306334
rect -5814 269778 -5258 270334
rect -5814 233778 -5258 234334
rect -5814 197778 -5258 198334
rect -5814 161778 -5258 162334
rect -5814 125778 -5258 126334
rect -5814 89778 -5258 90334
rect -5814 53778 -5258 54334
rect -5814 17778 -5258 18334
rect -4854 707162 -4298 707718
rect -4854 698058 -4298 698614
rect -4854 662058 -4298 662614
rect -4854 626058 -4298 626614
rect -4854 590058 -4298 590614
rect -4854 554058 -4298 554614
rect -4854 518058 -4298 518614
rect -4854 482058 -4298 482614
rect -4854 446058 -4298 446614
rect -4854 410058 -4298 410614
rect -4854 374058 -4298 374614
rect -4854 338058 -4298 338614
rect -4854 302058 -4298 302614
rect -4854 266058 -4298 266614
rect -4854 230058 -4298 230614
rect -4854 194058 -4298 194614
rect -4854 158058 -4298 158614
rect -4854 122058 -4298 122614
rect -4854 86058 -4298 86614
rect -4854 50058 -4298 50614
rect -4854 14058 -4298 14614
rect -3894 706202 -3338 706758
rect -3894 694338 -3338 694894
rect -3894 658338 -3338 658894
rect -3894 622338 -3338 622894
rect -3894 586338 -3338 586894
rect -3894 550338 -3338 550894
rect -3894 514338 -3338 514894
rect -3894 478338 -3338 478894
rect -3894 442338 -3338 442894
rect -3894 406338 -3338 406894
rect -3894 370338 -3338 370894
rect -3894 334338 -3338 334894
rect -3894 298338 -3338 298894
rect -3894 262338 -3338 262894
rect -3894 226338 -3338 226894
rect -3894 190338 -3338 190894
rect -3894 154338 -3338 154894
rect -3894 118338 -3338 118894
rect -3894 82338 -3338 82894
rect -3894 46338 -3338 46894
rect -3894 10338 -3338 10894
rect -2934 705242 -2378 705798
rect -2934 690618 -2378 691174
rect -2934 654618 -2378 655174
rect -2934 618618 -2378 619174
rect -2934 582618 -2378 583174
rect -2934 546618 -2378 547174
rect -2934 510618 -2378 511174
rect -2934 474618 -2378 475174
rect -2934 438618 -2378 439174
rect -2934 402618 -2378 403174
rect -2934 366618 -2378 367174
rect -2934 330618 -2378 331174
rect -2934 294618 -2378 295174
rect -2934 258618 -2378 259174
rect -2934 222618 -2378 223174
rect -2934 186618 -2378 187174
rect -2934 150618 -2378 151174
rect -2934 114618 -2378 115174
rect -2934 78618 -2378 79174
rect -2934 42618 -2378 43174
rect -2934 6618 -2378 7174
rect -1974 704282 -1418 704838
rect -1974 686898 -1418 687454
rect -1974 650898 -1418 651454
rect -1974 614898 -1418 615454
rect -1974 578898 -1418 579454
rect -1974 542898 -1418 543454
rect -1974 506898 -1418 507454
rect -1974 470898 -1418 471454
rect -1974 434898 -1418 435454
rect -1974 398898 -1418 399454
rect -1974 362898 -1418 363454
rect -1974 326898 -1418 327454
rect -1974 290898 -1418 291454
rect -1974 254898 -1418 255454
rect -1974 218898 -1418 219454
rect -1974 182898 -1418 183454
rect -1974 146898 -1418 147454
rect -1974 110898 -1418 111454
rect -1974 74898 -1418 75454
rect -1974 38898 -1418 39454
rect -1974 2898 -1418 3454
rect -1974 -902 -1418 -346
rect 1826 704282 2382 704838
rect 1826 686898 2382 687454
rect 1826 650898 2382 651454
rect 1826 614898 2382 615454
rect 1826 578898 2382 579454
rect 1826 542898 2382 543454
rect 1826 506898 2382 507454
rect 1826 470898 2382 471454
rect 1826 434898 2382 435454
rect 1826 398898 2382 399454
rect 1826 362898 2382 363454
rect 1826 326898 2382 327454
rect 1826 290898 2382 291454
rect 1826 254898 2382 255454
rect 1826 218898 2382 219454
rect 1826 182898 2382 183454
rect 1826 146898 2382 147454
rect 1826 110898 2382 111454
rect 1826 74898 2382 75454
rect 1826 38898 2382 39454
rect 1826 2898 2382 3454
rect 1826 -902 2382 -346
rect -2934 -1862 -2378 -1306
rect -3894 -2822 -3338 -2266
rect -4854 -3782 -4298 -3226
rect -5814 -4742 -5258 -4186
rect -6774 -5702 -6218 -5146
rect -7734 -6662 -7178 -6106
rect -8694 -7622 -8138 -7066
rect 5546 705242 6102 705798
rect 5546 690618 6102 691174
rect 5546 654618 6102 655174
rect 5546 618618 6102 619174
rect 5546 582618 6102 583174
rect 5546 546618 6102 547174
rect 5546 510618 6102 511174
rect 5546 474618 6102 475174
rect 5546 438618 6102 439174
rect 5546 402618 6102 403174
rect 5546 366618 6102 367174
rect 5546 330618 6102 331174
rect 5546 294618 6102 295174
rect 5546 258618 6102 259174
rect 5546 222618 6102 223174
rect 5546 186618 6102 187174
rect 5546 150618 6102 151174
rect 5546 114618 6102 115174
rect 5546 78618 6102 79174
rect 5546 42618 6102 43174
rect 5546 6618 6102 7174
rect 5546 -1862 6102 -1306
rect 9266 706202 9822 706758
rect 9266 694338 9822 694894
rect 9266 658338 9822 658894
rect 9266 622338 9822 622894
rect 9266 586338 9822 586894
rect 9266 550338 9822 550894
rect 9266 514338 9822 514894
rect 9266 478338 9822 478894
rect 9266 442338 9822 442894
rect 9266 406338 9822 406894
rect 9266 370338 9822 370894
rect 9266 334338 9822 334894
rect 9266 298338 9822 298894
rect 9266 262338 9822 262894
rect 9266 226338 9822 226894
rect 9266 190338 9822 190894
rect 9266 154338 9822 154894
rect 9266 118338 9822 118894
rect 9266 82338 9822 82894
rect 9266 46338 9822 46894
rect 9266 10338 9822 10894
rect 9266 -2822 9822 -2266
rect 12986 707162 13542 707718
rect 12986 698058 13542 698614
rect 12986 662058 13542 662614
rect 12986 626058 13542 626614
rect 12986 590058 13542 590614
rect 12986 554058 13542 554614
rect 12986 518058 13542 518614
rect 12986 482058 13542 482614
rect 12986 446058 13542 446614
rect 12986 410058 13542 410614
rect 12986 374058 13542 374614
rect 12986 338058 13542 338614
rect 12986 302058 13542 302614
rect 12986 266058 13542 266614
rect 16706 708122 17262 708678
rect 16706 665778 17262 666334
rect 16706 629778 17262 630334
rect 16706 593778 17262 594334
rect 16706 557778 17262 558334
rect 16706 521778 17262 522334
rect 16706 485778 17262 486334
rect 16706 449778 17262 450334
rect 16706 413778 17262 414334
rect 16706 377778 17262 378334
rect 16706 341778 17262 342334
rect 16706 305778 17262 306334
rect 16706 269778 17262 270334
rect 16250 255218 16486 255454
rect 16250 254898 16486 255134
rect 12986 230058 13542 230614
rect 16706 233778 17262 234334
rect 16250 219218 16486 219454
rect 16250 218898 16486 219134
rect 12986 194058 13542 194614
rect 16706 197778 17262 198334
rect 16250 183218 16486 183454
rect 16250 182898 16486 183134
rect 12986 158058 13542 158614
rect 16706 161778 17262 162334
rect 20426 709082 20982 709638
rect 20426 669498 20982 670054
rect 20426 633498 20982 634054
rect 20426 597498 20982 598054
rect 20426 561498 20982 562054
rect 20426 525498 20982 526054
rect 20426 489498 20982 490054
rect 20426 453498 20982 454054
rect 20426 417498 20982 418054
rect 20426 381498 20982 382054
rect 20426 345498 20982 346054
rect 20426 309498 20982 310054
rect 24146 710042 24702 710598
rect 24146 673218 24702 673774
rect 24146 637218 24702 637774
rect 24146 601218 24702 601774
rect 24146 565218 24702 565774
rect 24146 529218 24702 529774
rect 24146 493218 24702 493774
rect 24146 457218 24702 457774
rect 24146 421218 24702 421774
rect 24146 385218 24702 385774
rect 24146 349218 24702 349774
rect 24146 313218 24702 313774
rect 27866 711002 28422 711558
rect 27866 676938 28422 677494
rect 27866 640938 28422 641494
rect 27866 604938 28422 605494
rect 27866 568938 28422 569494
rect 27866 532938 28422 533494
rect 27866 496938 28422 497494
rect 27866 460938 28422 461494
rect 27866 424938 28422 425494
rect 27866 388938 28422 389494
rect 27866 352938 28422 353494
rect 27866 316938 28422 317494
rect 20426 273498 20982 274054
rect 27866 280938 28422 281494
rect 23930 258938 24166 259174
rect 23930 258618 24166 258854
rect 20426 237498 20982 238054
rect 37826 704282 38382 704838
rect 37826 686898 38382 687454
rect 37826 650898 38382 651454
rect 37826 614898 38382 615454
rect 37826 578898 38382 579454
rect 37826 542898 38382 543454
rect 37826 506898 38382 507454
rect 37826 470898 38382 471454
rect 37826 434898 38382 435454
rect 37826 398898 38382 399454
rect 37826 362898 38382 363454
rect 37826 326898 38382 327454
rect 37826 290898 38382 291454
rect 31610 270098 31846 270334
rect 31610 269778 31846 270014
rect 27866 244938 28422 245494
rect 23930 222938 24166 223174
rect 23930 222618 24166 222854
rect 20426 201498 20982 202054
rect 41546 705242 42102 705798
rect 41546 690618 42102 691174
rect 41546 654618 42102 655174
rect 41546 618618 42102 619174
rect 41546 582618 42102 583174
rect 41546 546618 42102 547174
rect 41546 510618 42102 511174
rect 41546 474618 42102 475174
rect 41546 438618 42102 439174
rect 41546 402618 42102 403174
rect 41546 366618 42102 367174
rect 41546 330618 42102 331174
rect 41546 294618 42102 295174
rect 39290 273818 39526 274054
rect 39290 273498 39526 273734
rect 37826 254898 38382 255454
rect 31610 234098 31846 234334
rect 31610 233778 31846 234014
rect 27866 208938 28422 209494
rect 23930 186938 24166 187174
rect 23930 186618 24166 186854
rect 20426 165498 20982 166054
rect 16250 147218 16486 147454
rect 16250 146898 16486 147134
rect 12986 122058 13542 122614
rect 41546 258618 42102 259174
rect 39290 237818 39526 238054
rect 39290 237498 39526 237734
rect 37826 218898 38382 219454
rect 31610 198098 31846 198334
rect 31610 197778 31846 198014
rect 27866 172938 28422 173494
rect 23930 150938 24166 151174
rect 23930 150618 24166 150854
rect 20426 129498 20982 130054
rect 17310 114938 17546 115174
rect 17310 114618 17546 114854
rect 16250 111218 16486 111454
rect 16250 110898 16486 111134
rect 12986 86058 13542 86614
rect 41546 222618 42102 223174
rect 39290 201818 39526 202054
rect 39290 201498 39526 201734
rect 37826 182898 38382 183454
rect 31610 162098 31846 162334
rect 31610 161778 31846 162014
rect 27866 136938 28422 137494
rect 23930 114938 24166 115174
rect 23930 114618 24166 114854
rect 20426 93498 20982 94054
rect 17310 78938 17546 79174
rect 17310 78618 17546 78854
rect 16250 75218 16486 75454
rect 16250 74898 16486 75134
rect 12986 50058 13542 50614
rect 41546 186618 42102 187174
rect 39290 165818 39526 166054
rect 39290 165498 39526 165734
rect 37826 146898 38382 147454
rect 31610 126098 31846 126334
rect 31610 125778 31846 126014
rect 27866 100938 28422 101494
rect 23930 78938 24166 79174
rect 23930 78618 24166 78854
rect 20426 57498 20982 58054
rect 17310 42938 17546 43174
rect 17310 42618 17546 42854
rect 16250 39218 16486 39454
rect 16250 38898 16486 39134
rect 12986 14058 13542 14614
rect 41546 150618 42102 151174
rect 39290 129818 39526 130054
rect 39290 129498 39526 129734
rect 37826 110898 38382 111454
rect 31610 90098 31846 90334
rect 31610 89778 31846 90014
rect 27866 64938 28422 65494
rect 23930 42938 24166 43174
rect 23930 42618 24166 42854
rect 20426 21498 20982 22054
rect 17310 6938 17546 7174
rect 17310 6618 17546 6854
rect 12986 -3782 13542 -3226
rect 16706 -4742 17262 -4186
rect 41546 114618 42102 115174
rect 39290 93818 39526 94054
rect 39290 93498 39526 93734
rect 37826 74898 38382 75454
rect 31610 54098 31846 54334
rect 31610 53778 31846 54014
rect 27866 28938 28422 29494
rect 23930 6938 24166 7174
rect 23930 6618 24166 6854
rect 20426 -5702 20982 -5146
rect 24146 -6662 24702 -6106
rect 41546 78618 42102 79174
rect 39290 57818 39526 58054
rect 39290 57498 39526 57734
rect 37826 38898 38382 39454
rect 31610 18098 31846 18334
rect 31610 17778 31846 18014
rect 27866 -7622 28422 -7066
rect 41546 42618 42102 43174
rect 39290 21818 39526 22054
rect 39290 21498 39526 21734
rect 37826 2898 38382 3454
rect 37826 -902 38382 -346
rect 41546 6618 42102 7174
rect 41546 -1862 42102 -1306
rect 45266 706202 45822 706758
rect 45266 694338 45822 694894
rect 45266 658338 45822 658894
rect 45266 622338 45822 622894
rect 45266 586338 45822 586894
rect 45266 550338 45822 550894
rect 45266 514338 45822 514894
rect 45266 478338 45822 478894
rect 45266 442338 45822 442894
rect 45266 406338 45822 406894
rect 45266 370338 45822 370894
rect 45266 334338 45822 334894
rect 45266 298338 45822 298894
rect 45266 262338 45822 262894
rect 48986 707162 49542 707718
rect 48986 698058 49542 698614
rect 48986 662058 49542 662614
rect 48986 626058 49542 626614
rect 48986 590058 49542 590614
rect 48986 554058 49542 554614
rect 48986 518058 49542 518614
rect 48986 482058 49542 482614
rect 48986 446058 49542 446614
rect 48986 410058 49542 410614
rect 48986 374058 49542 374614
rect 48986 338058 49542 338614
rect 48986 302058 49542 302614
rect 48986 266058 49542 266614
rect 46970 255218 47206 255454
rect 46970 254898 47206 255134
rect 45266 226338 45822 226894
rect 48986 230058 49542 230614
rect 46970 219218 47206 219454
rect 46970 218898 47206 219134
rect 45266 190338 45822 190894
rect 48986 194058 49542 194614
rect 46970 183218 47206 183454
rect 46970 182898 47206 183134
rect 45266 154338 45822 154894
rect 48986 158058 49542 158614
rect 46970 147218 47206 147454
rect 46970 146898 47206 147134
rect 45266 118338 45822 118894
rect 48986 122058 49542 122614
rect 46970 111218 47206 111454
rect 46970 110898 47206 111134
rect 45266 82338 45822 82894
rect 48986 86058 49542 86614
rect 46970 75218 47206 75454
rect 46970 74898 47206 75134
rect 45266 46338 45822 46894
rect 48986 50058 49542 50614
rect 46970 39218 47206 39454
rect 46970 38898 47206 39134
rect 45266 10338 45822 10894
rect 45266 -2822 45822 -2266
rect 48986 14058 49542 14614
rect 48986 -3782 49542 -3226
rect 52706 708122 53262 708678
rect 52706 665778 53262 666334
rect 52706 629778 53262 630334
rect 52706 593778 53262 594334
rect 52706 557778 53262 558334
rect 52706 521778 53262 522334
rect 52706 485778 53262 486334
rect 52706 449778 53262 450334
rect 52706 413778 53262 414334
rect 52706 377778 53262 378334
rect 52706 341778 53262 342334
rect 52706 305778 53262 306334
rect 52706 269778 53262 270334
rect 56426 709082 56982 709638
rect 56426 669498 56982 670054
rect 56426 633498 56982 634054
rect 56426 597498 56982 598054
rect 56426 561498 56982 562054
rect 56426 525498 56982 526054
rect 56426 489498 56982 490054
rect 56426 453498 56982 454054
rect 56426 417498 56982 418054
rect 56426 381498 56982 382054
rect 56426 345498 56982 346054
rect 56426 309498 56982 310054
rect 56426 273498 56982 274054
rect 54650 258938 54886 259174
rect 54650 258618 54886 258854
rect 52706 233778 53262 234334
rect 56426 237498 56982 238054
rect 54650 222938 54886 223174
rect 54650 222618 54886 222854
rect 52706 197778 53262 198334
rect 56426 201498 56982 202054
rect 54650 186938 54886 187174
rect 54650 186618 54886 186854
rect 52706 161778 53262 162334
rect 56426 165498 56982 166054
rect 54650 150938 54886 151174
rect 54650 150618 54886 150854
rect 52706 125778 53262 126334
rect 56426 129498 56982 130054
rect 54650 114938 54886 115174
rect 54650 114618 54886 114854
rect 52706 89778 53262 90334
rect 56426 93498 56982 94054
rect 54650 78938 54886 79174
rect 54650 78618 54886 78854
rect 52706 53778 53262 54334
rect 56426 57498 56982 58054
rect 54650 42938 54886 43174
rect 54650 42618 54886 42854
rect 52706 17778 53262 18334
rect 56426 21498 56982 22054
rect 54650 6938 54886 7174
rect 54650 6618 54886 6854
rect 52706 -4742 53262 -4186
rect 56426 -5702 56982 -5146
rect 60146 710042 60702 710598
rect 60146 673218 60702 673774
rect 60146 637218 60702 637774
rect 60146 601218 60702 601774
rect 60146 565218 60702 565774
rect 60146 529218 60702 529774
rect 60146 493218 60702 493774
rect 60146 457218 60702 457774
rect 60146 421218 60702 421774
rect 60146 385218 60702 385774
rect 60146 349218 60702 349774
rect 60146 313218 60702 313774
rect 60146 277218 60702 277774
rect 63866 711002 64422 711558
rect 63866 676938 64422 677494
rect 63866 640938 64422 641494
rect 63866 604938 64422 605494
rect 63866 568938 64422 569494
rect 63866 532938 64422 533494
rect 63866 496938 64422 497494
rect 63866 460938 64422 461494
rect 63866 424938 64422 425494
rect 63866 388938 64422 389494
rect 63866 352938 64422 353494
rect 63866 316938 64422 317494
rect 63866 280938 64422 281494
rect 62330 270098 62566 270334
rect 62330 269778 62566 270014
rect 60146 241218 60702 241774
rect 73826 704282 74382 704838
rect 73826 686898 74382 687454
rect 73826 650898 74382 651454
rect 73826 614898 74382 615454
rect 73826 578898 74382 579454
rect 73826 542898 74382 543454
rect 73826 506898 74382 507454
rect 73826 470898 74382 471454
rect 73826 434898 74382 435454
rect 73826 398898 74382 399454
rect 73826 362898 74382 363454
rect 73826 326898 74382 327454
rect 73826 290898 74382 291454
rect 70010 273818 70246 274054
rect 70010 273498 70246 273734
rect 63866 244938 64422 245494
rect 62330 234098 62566 234334
rect 62330 233778 62566 234014
rect 60146 205218 60702 205774
rect 77546 705242 78102 705798
rect 77546 690618 78102 691174
rect 77546 654618 78102 655174
rect 77546 618618 78102 619174
rect 77546 582618 78102 583174
rect 77546 546618 78102 547174
rect 77546 510618 78102 511174
rect 77546 474618 78102 475174
rect 77546 438618 78102 439174
rect 77546 402618 78102 403174
rect 77546 366618 78102 367174
rect 77546 330618 78102 331174
rect 77546 294618 78102 295174
rect 81266 706202 81822 706758
rect 81266 694338 81822 694894
rect 81266 658338 81822 658894
rect 81266 622338 81822 622894
rect 81266 586338 81822 586894
rect 81266 550338 81822 550894
rect 81266 514338 81822 514894
rect 81266 478338 81822 478894
rect 81266 442338 81822 442894
rect 81266 406338 81822 406894
rect 81266 370338 81822 370894
rect 81266 334338 81822 334894
rect 81266 298338 81822 298894
rect 84986 707162 85542 707718
rect 84986 698058 85542 698614
rect 84986 662058 85542 662614
rect 84986 626058 85542 626614
rect 84986 590058 85542 590614
rect 84986 554058 85542 554614
rect 84986 518058 85542 518614
rect 84986 482058 85542 482614
rect 84986 446058 85542 446614
rect 84986 410058 85542 410614
rect 84986 374058 85542 374614
rect 84986 338058 85542 338614
rect 84986 302058 85542 302614
rect 88706 708122 89262 708678
rect 88706 665778 89262 666334
rect 88706 629778 89262 630334
rect 88706 593778 89262 594334
rect 88706 557778 89262 558334
rect 88706 521778 89262 522334
rect 88706 485778 89262 486334
rect 88706 449778 89262 450334
rect 88706 413778 89262 414334
rect 88706 377778 89262 378334
rect 88706 341778 89262 342334
rect 88706 305778 89262 306334
rect 81266 262338 81822 262894
rect 73826 254898 74382 255454
rect 70010 237818 70246 238054
rect 70010 237498 70246 237734
rect 63866 208938 64422 209494
rect 62330 198098 62566 198334
rect 62330 197778 62566 198014
rect 60146 169218 60702 169774
rect 77690 255218 77926 255454
rect 77690 254898 77926 255134
rect 92426 709082 92982 709638
rect 92426 669498 92982 670054
rect 92426 633498 92982 634054
rect 92426 597498 92982 598054
rect 92426 561498 92982 562054
rect 92426 525498 92982 526054
rect 92426 489498 92982 490054
rect 92426 453498 92982 454054
rect 92426 417498 92982 418054
rect 92426 381498 92982 382054
rect 92426 345498 92982 346054
rect 92426 309498 92982 310054
rect 96146 710042 96702 710598
rect 96146 673218 96702 673774
rect 96146 637218 96702 637774
rect 96146 601218 96702 601774
rect 96146 565218 96702 565774
rect 96146 529218 96702 529774
rect 96146 493218 96702 493774
rect 96146 457218 96702 457774
rect 96146 421218 96702 421774
rect 96146 385218 96702 385774
rect 96146 349218 96702 349774
rect 96146 313218 96702 313774
rect 96146 277218 96702 277774
rect 88706 269778 89262 270334
rect 85370 258938 85606 259174
rect 85370 258618 85606 258854
rect 81266 226338 81822 226894
rect 73826 218898 74382 219454
rect 70010 201818 70246 202054
rect 70010 201498 70246 201734
rect 63866 172938 64422 173494
rect 62330 162098 62566 162334
rect 62330 161778 62566 162014
rect 60146 133218 60702 133774
rect 77690 219218 77926 219454
rect 77690 218898 77926 219134
rect 93050 270098 93286 270334
rect 93050 269778 93286 270014
rect 96146 241218 96702 241774
rect 88706 233778 89262 234334
rect 85370 222938 85606 223174
rect 85370 222618 85606 222854
rect 81266 190338 81822 190894
rect 73826 182898 74382 183454
rect 70010 165818 70246 166054
rect 70010 165498 70246 165734
rect 63866 136938 64422 137494
rect 62330 126098 62566 126334
rect 62330 125778 62566 126014
rect 60146 97218 60702 97774
rect 77690 183218 77926 183454
rect 77690 182898 77926 183134
rect 93050 234098 93286 234334
rect 93050 233778 93286 234014
rect 96146 205218 96702 205774
rect 88706 197778 89262 198334
rect 85370 186938 85606 187174
rect 85370 186618 85606 186854
rect 81266 154338 81822 154894
rect 73826 146898 74382 147454
rect 70010 129818 70246 130054
rect 70010 129498 70246 129734
rect 63866 100938 64422 101494
rect 62330 90098 62566 90334
rect 62330 89778 62566 90014
rect 60146 61218 60702 61774
rect 77690 147218 77926 147454
rect 77690 146898 77926 147134
rect 93050 198098 93286 198334
rect 93050 197778 93286 198014
rect 96146 169218 96702 169774
rect 88706 161778 89262 162334
rect 85370 150938 85606 151174
rect 85370 150618 85606 150854
rect 81266 118338 81822 118894
rect 73826 110898 74382 111454
rect 70010 93818 70246 94054
rect 70010 93498 70246 93734
rect 63866 64938 64422 65494
rect 62330 54098 62566 54334
rect 62330 53778 62566 54014
rect 60146 25218 60702 25774
rect 77690 111218 77926 111454
rect 77690 110898 77926 111134
rect 93050 162098 93286 162334
rect 93050 161778 93286 162014
rect 96146 133218 96702 133774
rect 88706 125778 89262 126334
rect 85370 114938 85606 115174
rect 85370 114618 85606 114854
rect 81266 82338 81822 82894
rect 73826 74898 74382 75454
rect 70010 57818 70246 58054
rect 70010 57498 70246 57734
rect 63866 28938 64422 29494
rect 62330 18098 62566 18334
rect 62330 17778 62566 18014
rect 60146 -6662 60702 -6106
rect 77690 75218 77926 75454
rect 77690 74898 77926 75134
rect 93050 126098 93286 126334
rect 93050 125778 93286 126014
rect 96146 97218 96702 97774
rect 88706 89778 89262 90334
rect 85370 78938 85606 79174
rect 85370 78618 85606 78854
rect 81266 46338 81822 46894
rect 73826 38898 74382 39454
rect 70010 21818 70246 22054
rect 70010 21498 70246 21734
rect 63866 -7622 64422 -7066
rect 77690 39218 77926 39454
rect 77690 38898 77926 39134
rect 73826 2898 74382 3454
rect 93050 90098 93286 90334
rect 93050 89778 93286 90014
rect 96146 61218 96702 61774
rect 88706 53778 89262 54334
rect 85370 42938 85606 43174
rect 85370 42618 85606 42854
rect 81266 10338 81822 10894
rect 73826 -902 74382 -346
rect 77546 -1862 78102 -1306
rect 93050 54098 93286 54334
rect 93050 53778 93286 54014
rect 96146 25218 96702 25774
rect 88706 17778 89262 18334
rect 85370 6938 85606 7174
rect 85370 6618 85606 6854
rect 81266 -2822 81822 -2266
rect 84986 -3782 85542 -3226
rect 93050 18098 93286 18334
rect 93050 17778 93286 18014
rect 88706 -4742 89262 -4186
rect 92426 -5702 92982 -5146
rect 96146 -6662 96702 -6106
rect 99866 711002 100422 711558
rect 99866 676938 100422 677494
rect 99866 640938 100422 641494
rect 99866 604938 100422 605494
rect 99866 568938 100422 569494
rect 99866 532938 100422 533494
rect 99866 496938 100422 497494
rect 99866 460938 100422 461494
rect 99866 424938 100422 425494
rect 99866 388938 100422 389494
rect 99866 352938 100422 353494
rect 99866 316938 100422 317494
rect 99866 280938 100422 281494
rect 109826 704282 110382 704838
rect 109826 686898 110382 687454
rect 109826 650898 110382 651454
rect 109826 614898 110382 615454
rect 109826 578898 110382 579454
rect 109826 542898 110382 543454
rect 109826 506898 110382 507454
rect 109826 470898 110382 471454
rect 109826 434898 110382 435454
rect 109826 398898 110382 399454
rect 109826 362898 110382 363454
rect 109826 326898 110382 327454
rect 109826 290898 110382 291454
rect 100730 273818 100966 274054
rect 100730 273498 100966 273734
rect 108410 255218 108646 255454
rect 108410 254898 108646 255134
rect 109826 254898 110382 255454
rect 99866 244938 100422 245494
rect 100730 237818 100966 238054
rect 100730 237498 100966 237734
rect 108410 219218 108646 219454
rect 108410 218898 108646 219134
rect 109826 218898 110382 219454
rect 99866 208938 100422 209494
rect 100730 201818 100966 202054
rect 100730 201498 100966 201734
rect 108410 183218 108646 183454
rect 108410 182898 108646 183134
rect 109826 182898 110382 183454
rect 99866 172938 100422 173494
rect 100730 165818 100966 166054
rect 100730 165498 100966 165734
rect 108410 147218 108646 147454
rect 108410 146898 108646 147134
rect 109826 146898 110382 147454
rect 99866 136938 100422 137494
rect 100730 129818 100966 130054
rect 100730 129498 100966 129734
rect 108410 111218 108646 111454
rect 108410 110898 108646 111134
rect 113546 705242 114102 705798
rect 113546 690618 114102 691174
rect 113546 654618 114102 655174
rect 113546 618618 114102 619174
rect 113546 582618 114102 583174
rect 113546 546618 114102 547174
rect 113546 510618 114102 511174
rect 113546 474618 114102 475174
rect 113546 438618 114102 439174
rect 113546 402618 114102 403174
rect 113546 366618 114102 367174
rect 113546 330618 114102 331174
rect 113546 294618 114102 295174
rect 117266 706202 117822 706758
rect 117266 694338 117822 694894
rect 117266 658338 117822 658894
rect 117266 622338 117822 622894
rect 117266 586338 117822 586894
rect 117266 550338 117822 550894
rect 117266 514338 117822 514894
rect 117266 478338 117822 478894
rect 117266 442338 117822 442894
rect 117266 406338 117822 406894
rect 117266 370338 117822 370894
rect 117266 334338 117822 334894
rect 117266 298338 117822 298894
rect 117266 262338 117822 262894
rect 113546 258618 114102 259174
rect 116090 258938 116326 259174
rect 116090 258618 116326 258854
rect 117266 226338 117822 226894
rect 113546 222618 114102 223174
rect 116090 222938 116326 223174
rect 116090 222618 116326 222854
rect 117266 190338 117822 190894
rect 113546 186618 114102 187174
rect 116090 186938 116326 187174
rect 116090 186618 116326 186854
rect 117266 154338 117822 154894
rect 113546 150618 114102 151174
rect 116090 150938 116326 151174
rect 116090 150618 116326 150854
rect 117266 118338 117822 118894
rect 116090 114938 116326 115174
rect 116090 114618 116326 114854
rect 109826 110898 110382 111454
rect 99866 100938 100422 101494
rect 100730 93818 100966 94054
rect 100730 93498 100966 93734
rect 108410 75218 108646 75454
rect 108410 74898 108646 75134
rect 117266 82338 117822 82894
rect 116090 78938 116326 79174
rect 116090 78618 116326 78854
rect 109826 74898 110382 75454
rect 99866 64938 100422 65494
rect 100730 57818 100966 58054
rect 100730 57498 100966 57734
rect 108410 39218 108646 39454
rect 108410 38898 108646 39134
rect 117266 46338 117822 46894
rect 116090 42938 116326 43174
rect 116090 42618 116326 42854
rect 109826 38898 110382 39454
rect 99866 28938 100422 29494
rect 100730 21818 100966 22054
rect 100730 21498 100966 21734
rect 99866 -7622 100422 -7066
rect 117266 10338 117822 10894
rect 116090 6938 116326 7174
rect 116090 6618 116326 6854
rect 109826 2898 110382 3454
rect 109826 -902 110382 -346
rect 113546 -1862 114102 -1306
rect 117266 -2822 117822 -2266
rect 120986 707162 121542 707718
rect 120986 698058 121542 698614
rect 120986 662058 121542 662614
rect 120986 626058 121542 626614
rect 120986 590058 121542 590614
rect 120986 554058 121542 554614
rect 120986 518058 121542 518614
rect 120986 482058 121542 482614
rect 120986 446058 121542 446614
rect 120986 410058 121542 410614
rect 120986 374058 121542 374614
rect 120986 338058 121542 338614
rect 120986 302058 121542 302614
rect 124706 708122 125262 708678
rect 124706 665778 125262 666334
rect 124706 629778 125262 630334
rect 124706 593778 125262 594334
rect 124706 557778 125262 558334
rect 124706 521778 125262 522334
rect 124706 485778 125262 486334
rect 124706 449778 125262 450334
rect 124706 413778 125262 414334
rect 124706 377778 125262 378334
rect 124706 341778 125262 342334
rect 124706 305778 125262 306334
rect 123770 270098 124006 270334
rect 123770 269778 124006 270014
rect 124706 269778 125262 270334
rect 120986 266058 121542 266614
rect 123770 234098 124006 234334
rect 123770 233778 124006 234014
rect 124706 233778 125262 234334
rect 120986 230058 121542 230614
rect 123770 198098 124006 198334
rect 123770 197778 124006 198014
rect 124706 197778 125262 198334
rect 120986 194058 121542 194614
rect 123770 162098 124006 162334
rect 123770 161778 124006 162014
rect 124706 161778 125262 162334
rect 120986 158058 121542 158614
rect 123770 126098 124006 126334
rect 123770 125778 124006 126014
rect 124706 125778 125262 126334
rect 120986 122058 121542 122614
rect 123770 90098 124006 90334
rect 123770 89778 124006 90014
rect 124706 89778 125262 90334
rect 120986 86058 121542 86614
rect 123770 54098 124006 54334
rect 123770 53778 124006 54014
rect 124706 53778 125262 54334
rect 120986 50058 121542 50614
rect 123770 18098 124006 18334
rect 123770 17778 124006 18014
rect 124706 17778 125262 18334
rect 120986 14058 121542 14614
rect 120986 -3782 121542 -3226
rect 124706 -4742 125262 -4186
rect 128426 709082 128982 709638
rect 128426 669498 128982 670054
rect 128426 633498 128982 634054
rect 128426 597498 128982 598054
rect 128426 561498 128982 562054
rect 128426 525498 128982 526054
rect 128426 489498 128982 490054
rect 128426 453498 128982 454054
rect 128426 417498 128982 418054
rect 128426 381498 128982 382054
rect 128426 345498 128982 346054
rect 128426 309498 128982 310054
rect 132146 710042 132702 710598
rect 132146 673218 132702 673774
rect 132146 637218 132702 637774
rect 132146 601218 132702 601774
rect 132146 565218 132702 565774
rect 132146 529218 132702 529774
rect 132146 493218 132702 493774
rect 132146 457218 132702 457774
rect 132146 421218 132702 421774
rect 132146 385218 132702 385774
rect 132146 349218 132702 349774
rect 132146 313218 132702 313774
rect 132146 277218 132702 277774
rect 128426 273498 128982 274054
rect 131450 273818 131686 274054
rect 131450 273498 131686 273734
rect 132146 241218 132702 241774
rect 128426 237498 128982 238054
rect 131450 237818 131686 238054
rect 131450 237498 131686 237734
rect 132146 205218 132702 205774
rect 128426 201498 128982 202054
rect 131450 201818 131686 202054
rect 131450 201498 131686 201734
rect 132146 169218 132702 169774
rect 128426 165498 128982 166054
rect 131450 165818 131686 166054
rect 131450 165498 131686 165734
rect 132146 133218 132702 133774
rect 128426 129498 128982 130054
rect 131450 129818 131686 130054
rect 131450 129498 131686 129734
rect 132146 97218 132702 97774
rect 128426 93498 128982 94054
rect 131450 93818 131686 94054
rect 131450 93498 131686 93734
rect 132146 61218 132702 61774
rect 128426 57498 128982 58054
rect 131450 57818 131686 58054
rect 131450 57498 131686 57734
rect 132146 25218 132702 25774
rect 128426 21498 128982 22054
rect 131450 21818 131686 22054
rect 131450 21498 131686 21734
rect 128426 -5702 128982 -5146
rect 132146 -6662 132702 -6106
rect 135866 711002 136422 711558
rect 135866 676938 136422 677494
rect 135866 640938 136422 641494
rect 135866 604938 136422 605494
rect 135866 568938 136422 569494
rect 135866 532938 136422 533494
rect 135866 496938 136422 497494
rect 135866 460938 136422 461494
rect 135866 424938 136422 425494
rect 135866 388938 136422 389494
rect 135866 352938 136422 353494
rect 135866 316938 136422 317494
rect 135866 280938 136422 281494
rect 145826 704282 146382 704838
rect 145826 686898 146382 687454
rect 145826 650898 146382 651454
rect 145826 614898 146382 615454
rect 145826 578898 146382 579454
rect 145826 542898 146382 543454
rect 145826 506898 146382 507454
rect 145826 470898 146382 471454
rect 145826 434898 146382 435454
rect 145826 398898 146382 399454
rect 145826 362898 146382 363454
rect 145826 326898 146382 327454
rect 145826 290898 146382 291454
rect 139130 255218 139366 255454
rect 139130 254898 139366 255134
rect 149546 705242 150102 705798
rect 149546 690618 150102 691174
rect 149546 654618 150102 655174
rect 149546 618618 150102 619174
rect 149546 582618 150102 583174
rect 149546 546618 150102 547174
rect 149546 510618 150102 511174
rect 149546 474618 150102 475174
rect 149546 438618 150102 439174
rect 149546 402618 150102 403174
rect 149546 366618 150102 367174
rect 149546 330618 150102 331174
rect 149546 294618 150102 295174
rect 146810 258938 147046 259174
rect 146810 258618 147046 258854
rect 149546 258618 150102 259174
rect 145826 254898 146382 255454
rect 135866 244938 136422 245494
rect 139130 219218 139366 219454
rect 139130 218898 139366 219134
rect 146810 222938 147046 223174
rect 146810 222618 147046 222854
rect 149546 222618 150102 223174
rect 145826 218898 146382 219454
rect 135866 208938 136422 209494
rect 139130 183218 139366 183454
rect 139130 182898 139366 183134
rect 146810 186938 147046 187174
rect 146810 186618 147046 186854
rect 149546 186618 150102 187174
rect 145826 182898 146382 183454
rect 135866 172938 136422 173494
rect 139130 147218 139366 147454
rect 139130 146898 139366 147134
rect 146810 150938 147046 151174
rect 146810 150618 147046 150854
rect 149546 150618 150102 151174
rect 145826 146898 146382 147454
rect 135866 136938 136422 137494
rect 139130 111218 139366 111454
rect 139130 110898 139366 111134
rect 146810 114938 147046 115174
rect 146810 114618 147046 114854
rect 149546 114618 150102 115174
rect 145826 110898 146382 111454
rect 135866 100938 136422 101494
rect 139130 75218 139366 75454
rect 139130 74898 139366 75134
rect 146810 78938 147046 79174
rect 146810 78618 147046 78854
rect 149546 78618 150102 79174
rect 145826 74898 146382 75454
rect 135866 64938 136422 65494
rect 139130 39218 139366 39454
rect 139130 38898 139366 39134
rect 146810 42938 147046 43174
rect 146810 42618 147046 42854
rect 149546 42618 150102 43174
rect 145826 38898 146382 39454
rect 135866 28938 136422 29494
rect 135866 -7622 136422 -7066
rect 146810 6938 147046 7174
rect 146810 6618 147046 6854
rect 149546 6618 150102 7174
rect 145826 2898 146382 3454
rect 145826 -902 146382 -346
rect 149546 -1862 150102 -1306
rect 153266 706202 153822 706758
rect 153266 694338 153822 694894
rect 153266 658338 153822 658894
rect 153266 622338 153822 622894
rect 153266 586338 153822 586894
rect 153266 550338 153822 550894
rect 153266 514338 153822 514894
rect 153266 478338 153822 478894
rect 153266 442338 153822 442894
rect 153266 406338 153822 406894
rect 153266 370338 153822 370894
rect 153266 334338 153822 334894
rect 153266 298338 153822 298894
rect 156986 707162 157542 707718
rect 156986 698058 157542 698614
rect 156986 662058 157542 662614
rect 156986 626058 157542 626614
rect 156986 590058 157542 590614
rect 156986 554058 157542 554614
rect 156986 518058 157542 518614
rect 156986 482058 157542 482614
rect 156986 446058 157542 446614
rect 156986 410058 157542 410614
rect 156986 374058 157542 374614
rect 156986 338058 157542 338614
rect 156986 302058 157542 302614
rect 154490 270098 154726 270334
rect 154490 269778 154726 270014
rect 153266 262338 153822 262894
rect 156986 266058 157542 266614
rect 154490 234098 154726 234334
rect 154490 233778 154726 234014
rect 153266 226338 153822 226894
rect 156986 230058 157542 230614
rect 154490 198098 154726 198334
rect 154490 197778 154726 198014
rect 153266 190338 153822 190894
rect 156986 194058 157542 194614
rect 154490 162098 154726 162334
rect 154490 161778 154726 162014
rect 153266 154338 153822 154894
rect 156986 158058 157542 158614
rect 154490 126098 154726 126334
rect 154490 125778 154726 126014
rect 153266 118338 153822 118894
rect 156986 122058 157542 122614
rect 154490 90098 154726 90334
rect 154490 89778 154726 90014
rect 153266 82338 153822 82894
rect 156986 86058 157542 86614
rect 154490 54098 154726 54334
rect 154490 53778 154726 54014
rect 153266 46338 153822 46894
rect 156986 50058 157542 50614
rect 154490 18098 154726 18334
rect 154490 17778 154726 18014
rect 153266 10338 153822 10894
rect 153266 -2822 153822 -2266
rect 156986 14058 157542 14614
rect 156986 -3782 157542 -3226
rect 160706 708122 161262 708678
rect 160706 665778 161262 666334
rect 160706 629778 161262 630334
rect 160706 593778 161262 594334
rect 160706 557778 161262 558334
rect 160706 521778 161262 522334
rect 160706 485778 161262 486334
rect 160706 449778 161262 450334
rect 160706 413778 161262 414334
rect 160706 377778 161262 378334
rect 160706 341778 161262 342334
rect 160706 305778 161262 306334
rect 164426 709082 164982 709638
rect 164426 669498 164982 670054
rect 164426 633498 164982 634054
rect 164426 597498 164982 598054
rect 164426 561498 164982 562054
rect 164426 525498 164982 526054
rect 164426 489498 164982 490054
rect 164426 453498 164982 454054
rect 164426 417498 164982 418054
rect 164426 381498 164982 382054
rect 164426 345498 164982 346054
rect 164426 309498 164982 310054
rect 162170 273818 162406 274054
rect 162170 273498 162406 273734
rect 164426 273498 164982 274054
rect 160706 269778 161262 270334
rect 162170 237818 162406 238054
rect 162170 237498 162406 237734
rect 164426 237498 164982 238054
rect 160706 233778 161262 234334
rect 162170 201818 162406 202054
rect 162170 201498 162406 201734
rect 164426 201498 164982 202054
rect 160706 197778 161262 198334
rect 162170 165818 162406 166054
rect 162170 165498 162406 165734
rect 164426 165498 164982 166054
rect 160706 161778 161262 162334
rect 162170 129818 162406 130054
rect 162170 129498 162406 129734
rect 164426 129498 164982 130054
rect 160706 125778 161262 126334
rect 162170 93818 162406 94054
rect 162170 93498 162406 93734
rect 164426 93498 164982 94054
rect 160706 89778 161262 90334
rect 162170 57818 162406 58054
rect 162170 57498 162406 57734
rect 164426 57498 164982 58054
rect 160706 53778 161262 54334
rect 162170 21818 162406 22054
rect 162170 21498 162406 21734
rect 164426 21498 164982 22054
rect 160706 17778 161262 18334
rect 160706 -4742 161262 -4186
rect 164426 -5702 164982 -5146
rect 168146 710042 168702 710598
rect 168146 673218 168702 673774
rect 168146 637218 168702 637774
rect 168146 601218 168702 601774
rect 168146 565218 168702 565774
rect 168146 529218 168702 529774
rect 168146 493218 168702 493774
rect 168146 457218 168702 457774
rect 168146 421218 168702 421774
rect 168146 385218 168702 385774
rect 168146 349218 168702 349774
rect 168146 313218 168702 313774
rect 168146 277218 168702 277774
rect 171866 711002 172422 711558
rect 171866 676938 172422 677494
rect 171866 640938 172422 641494
rect 171866 604938 172422 605494
rect 171866 568938 172422 569494
rect 171866 532938 172422 533494
rect 171866 496938 172422 497494
rect 171866 460938 172422 461494
rect 171866 424938 172422 425494
rect 171866 388938 172422 389494
rect 171866 352938 172422 353494
rect 171866 316938 172422 317494
rect 171866 280938 172422 281494
rect 169850 255218 170086 255454
rect 169850 254898 170086 255134
rect 168146 241218 168702 241774
rect 181826 704282 182382 704838
rect 181826 686898 182382 687454
rect 181826 650898 182382 651454
rect 181826 614898 182382 615454
rect 181826 578898 182382 579454
rect 181826 542898 182382 543454
rect 181826 506898 182382 507454
rect 181826 470898 182382 471454
rect 181826 434898 182382 435454
rect 181826 398898 182382 399454
rect 181826 362898 182382 363454
rect 181826 326898 182382 327454
rect 181826 290898 182382 291454
rect 177530 258938 177766 259174
rect 177530 258618 177766 258854
rect 171866 244938 172422 245494
rect 169850 219218 170086 219454
rect 169850 218898 170086 219134
rect 168146 205218 168702 205774
rect 185546 705242 186102 705798
rect 185546 690618 186102 691174
rect 185546 654618 186102 655174
rect 185546 618618 186102 619174
rect 185546 582618 186102 583174
rect 185546 546618 186102 547174
rect 185546 510618 186102 511174
rect 185546 474618 186102 475174
rect 185546 438618 186102 439174
rect 185546 402618 186102 403174
rect 185546 366618 186102 367174
rect 185546 330618 186102 331174
rect 185546 294618 186102 295174
rect 189266 706202 189822 706758
rect 189266 694338 189822 694894
rect 189266 658338 189822 658894
rect 189266 622338 189822 622894
rect 189266 586338 189822 586894
rect 189266 550338 189822 550894
rect 189266 514338 189822 514894
rect 189266 478338 189822 478894
rect 189266 442338 189822 442894
rect 189266 406338 189822 406894
rect 189266 370338 189822 370894
rect 189266 334338 189822 334894
rect 189266 298338 189822 298894
rect 185210 270098 185446 270334
rect 185210 269778 185446 270014
rect 181826 254898 182382 255454
rect 177530 222938 177766 223174
rect 177530 222618 177766 222854
rect 171866 208938 172422 209494
rect 169850 183218 170086 183454
rect 169850 182898 170086 183134
rect 168146 169218 168702 169774
rect 192986 707162 193542 707718
rect 192986 698058 193542 698614
rect 192986 662058 193542 662614
rect 192986 626058 193542 626614
rect 192986 590058 193542 590614
rect 192986 554058 193542 554614
rect 192986 518058 193542 518614
rect 192986 482058 193542 482614
rect 192986 446058 193542 446614
rect 192986 410058 193542 410614
rect 192986 374058 193542 374614
rect 192986 338058 193542 338614
rect 192986 302058 193542 302614
rect 196706 708122 197262 708678
rect 196706 665778 197262 666334
rect 196706 629778 197262 630334
rect 196706 593778 197262 594334
rect 196706 557778 197262 558334
rect 196706 521778 197262 522334
rect 196706 485778 197262 486334
rect 196706 449778 197262 450334
rect 196706 413778 197262 414334
rect 196706 377778 197262 378334
rect 196706 341778 197262 342334
rect 196706 305778 197262 306334
rect 192890 273818 193126 274054
rect 192890 273498 193126 273734
rect 189266 262338 189822 262894
rect 185210 234098 185446 234334
rect 185210 233778 185446 234014
rect 181826 218898 182382 219454
rect 177530 186938 177766 187174
rect 177530 186618 177766 186854
rect 171866 172938 172422 173494
rect 169850 147218 170086 147454
rect 169850 146898 170086 147134
rect 168146 133218 168702 133774
rect 200426 709082 200982 709638
rect 200426 669498 200982 670054
rect 200426 633498 200982 634054
rect 200426 597498 200982 598054
rect 200426 561498 200982 562054
rect 200426 525498 200982 526054
rect 200426 489498 200982 490054
rect 200426 453498 200982 454054
rect 200426 417498 200982 418054
rect 200426 381498 200982 382054
rect 200426 345498 200982 346054
rect 200426 309498 200982 310054
rect 204146 710042 204702 710598
rect 204146 673218 204702 673774
rect 204146 637218 204702 637774
rect 204146 601218 204702 601774
rect 204146 565218 204702 565774
rect 204146 529218 204702 529774
rect 204146 493218 204702 493774
rect 204146 457218 204702 457774
rect 204146 421218 204702 421774
rect 204146 385218 204702 385774
rect 204146 349218 204702 349774
rect 204146 313218 204702 313774
rect 196706 269778 197262 270334
rect 192890 237818 193126 238054
rect 192890 237498 193126 237734
rect 189266 226338 189822 226894
rect 185210 198098 185446 198334
rect 185210 197778 185446 198014
rect 181826 182898 182382 183454
rect 177530 150938 177766 151174
rect 177530 150618 177766 150854
rect 171866 136938 172422 137494
rect 169850 111218 170086 111454
rect 169850 110898 170086 111134
rect 168146 97218 168702 97774
rect 207866 711002 208422 711558
rect 207866 676938 208422 677494
rect 207866 640938 208422 641494
rect 207866 604938 208422 605494
rect 207866 568938 208422 569494
rect 207866 532938 208422 533494
rect 207866 496938 208422 497494
rect 207866 460938 208422 461494
rect 207866 424938 208422 425494
rect 207866 388938 208422 389494
rect 207866 352938 208422 353494
rect 207866 316938 208422 317494
rect 217826 704282 218382 704838
rect 217826 686898 218382 687454
rect 217826 650898 218382 651454
rect 217826 614898 218382 615454
rect 217826 578898 218382 579454
rect 217826 542898 218382 543454
rect 217826 506898 218382 507454
rect 217826 470898 218382 471454
rect 217826 434898 218382 435454
rect 217826 398898 218382 399454
rect 217826 362898 218382 363454
rect 217826 326898 218382 327454
rect 217826 290898 218382 291454
rect 204146 277218 204702 277774
rect 200570 255218 200806 255454
rect 200570 254898 200806 255134
rect 196706 233778 197262 234334
rect 192890 201818 193126 202054
rect 192890 201498 193126 201734
rect 189266 190338 189822 190894
rect 185210 162098 185446 162334
rect 185210 161778 185446 162014
rect 181826 146898 182382 147454
rect 177530 114938 177766 115174
rect 177530 114618 177766 114854
rect 171866 100938 172422 101494
rect 169850 75218 170086 75454
rect 169850 74898 170086 75134
rect 168146 61218 168702 61774
rect 215930 270098 216166 270334
rect 215930 269778 216166 270014
rect 208250 258938 208486 259174
rect 208250 258618 208486 258854
rect 204146 241218 204702 241774
rect 200570 219218 200806 219454
rect 200570 218898 200806 219134
rect 196706 197778 197262 198334
rect 192890 165818 193126 166054
rect 192890 165498 193126 165734
rect 189266 154338 189822 154894
rect 185210 126098 185446 126334
rect 185210 125778 185446 126014
rect 181826 110898 182382 111454
rect 177530 78938 177766 79174
rect 177530 78618 177766 78854
rect 171866 64938 172422 65494
rect 169850 39218 170086 39454
rect 169850 38898 170086 39134
rect 168146 25218 168702 25774
rect 168146 -6662 168702 -6106
rect 217826 254898 218382 255454
rect 215930 234098 216166 234334
rect 215930 233778 216166 234014
rect 208250 222938 208486 223174
rect 208250 222618 208486 222854
rect 204146 205218 204702 205774
rect 200570 183218 200806 183454
rect 200570 182898 200806 183134
rect 196706 161778 197262 162334
rect 192890 129818 193126 130054
rect 192890 129498 193126 129734
rect 189266 118338 189822 118894
rect 185210 90098 185446 90334
rect 185210 89778 185446 90014
rect 181826 74898 182382 75454
rect 177530 42938 177766 43174
rect 177530 42618 177766 42854
rect 171866 28938 172422 29494
rect 217826 218898 218382 219454
rect 215930 198098 216166 198334
rect 215930 197778 216166 198014
rect 208250 186938 208486 187174
rect 208250 186618 208486 186854
rect 204146 169218 204702 169774
rect 200570 147218 200806 147454
rect 200570 146898 200806 147134
rect 196706 125778 197262 126334
rect 192890 93818 193126 94054
rect 192890 93498 193126 93734
rect 189266 82338 189822 82894
rect 185210 54098 185446 54334
rect 185210 53778 185446 54014
rect 181826 38898 182382 39454
rect 177530 6938 177766 7174
rect 177530 6618 177766 6854
rect 171866 -7622 172422 -7066
rect 217826 182898 218382 183454
rect 215930 162098 216166 162334
rect 215930 161778 216166 162014
rect 208250 150938 208486 151174
rect 208250 150618 208486 150854
rect 204146 133218 204702 133774
rect 200570 111218 200806 111454
rect 200570 110898 200806 111134
rect 196706 89778 197262 90334
rect 192890 57818 193126 58054
rect 192890 57498 193126 57734
rect 189266 46338 189822 46894
rect 185210 18098 185446 18334
rect 185210 17778 185446 18014
rect 181826 2898 182382 3454
rect 217826 146898 218382 147454
rect 215930 126098 216166 126334
rect 215930 125778 216166 126014
rect 208250 114938 208486 115174
rect 208250 114618 208486 114854
rect 204146 97218 204702 97774
rect 200570 75218 200806 75454
rect 200570 74898 200806 75134
rect 196706 53778 197262 54334
rect 192890 21818 193126 22054
rect 192890 21498 193126 21734
rect 189266 10338 189822 10894
rect 181826 -902 182382 -346
rect 185546 -1862 186102 -1306
rect 217826 110898 218382 111454
rect 215930 90098 216166 90334
rect 215930 89778 216166 90014
rect 208250 78938 208486 79174
rect 208250 78618 208486 78854
rect 204146 61218 204702 61774
rect 200570 39218 200806 39454
rect 200570 38898 200806 39134
rect 196706 17778 197262 18334
rect 189266 -2822 189822 -2266
rect 192986 -3782 193542 -3226
rect 217826 74898 218382 75454
rect 215930 54098 216166 54334
rect 215930 53778 216166 54014
rect 208250 42938 208486 43174
rect 208250 42618 208486 42854
rect 204146 25218 204702 25774
rect 196706 -4742 197262 -4186
rect 200426 -5702 200982 -5146
rect 217826 38898 218382 39454
rect 215930 18098 216166 18334
rect 215930 17778 216166 18014
rect 208250 6938 208486 7174
rect 208250 6618 208486 6854
rect 204146 -6662 204702 -6106
rect 207866 -7622 208422 -7066
rect 217826 2898 218382 3454
rect 217826 -902 218382 -346
rect 221546 705242 222102 705798
rect 221546 690618 222102 691174
rect 221546 654618 222102 655174
rect 221546 618618 222102 619174
rect 221546 582618 222102 583174
rect 221546 546618 222102 547174
rect 221546 510618 222102 511174
rect 221546 474618 222102 475174
rect 221546 438618 222102 439174
rect 221546 402618 222102 403174
rect 221546 366618 222102 367174
rect 221546 330618 222102 331174
rect 221546 294618 222102 295174
rect 225266 706202 225822 706758
rect 225266 694338 225822 694894
rect 225266 658338 225822 658894
rect 225266 622338 225822 622894
rect 225266 586338 225822 586894
rect 225266 550338 225822 550894
rect 225266 514338 225822 514894
rect 225266 478338 225822 478894
rect 225266 442338 225822 442894
rect 225266 406338 225822 406894
rect 225266 370338 225822 370894
rect 225266 334338 225822 334894
rect 225266 298338 225822 298894
rect 223610 273818 223846 274054
rect 223610 273498 223846 273734
rect 221546 258618 222102 259174
rect 225266 262338 225822 262894
rect 223610 237818 223846 238054
rect 223610 237498 223846 237734
rect 221546 222618 222102 223174
rect 225266 226338 225822 226894
rect 223610 201818 223846 202054
rect 223610 201498 223846 201734
rect 221546 186618 222102 187174
rect 225266 190338 225822 190894
rect 223610 165818 223846 166054
rect 223610 165498 223846 165734
rect 221546 150618 222102 151174
rect 225266 154338 225822 154894
rect 223610 129818 223846 130054
rect 223610 129498 223846 129734
rect 221546 114618 222102 115174
rect 225266 118338 225822 118894
rect 223610 93818 223846 94054
rect 223610 93498 223846 93734
rect 221546 78618 222102 79174
rect 225266 82338 225822 82894
rect 223610 57818 223846 58054
rect 223610 57498 223846 57734
rect 221546 42618 222102 43174
rect 225266 46338 225822 46894
rect 223610 21818 223846 22054
rect 223610 21498 223846 21734
rect 221546 6618 222102 7174
rect 221546 -1862 222102 -1306
rect 225266 10338 225822 10894
rect 225266 -2822 225822 -2266
rect 228986 707162 229542 707718
rect 228986 698058 229542 698614
rect 228986 662058 229542 662614
rect 228986 626058 229542 626614
rect 228986 590058 229542 590614
rect 228986 554058 229542 554614
rect 228986 518058 229542 518614
rect 228986 482058 229542 482614
rect 228986 446058 229542 446614
rect 228986 410058 229542 410614
rect 228986 374058 229542 374614
rect 228986 338058 229542 338614
rect 228986 302058 229542 302614
rect 228986 266058 229542 266614
rect 232706 708122 233262 708678
rect 232706 665778 233262 666334
rect 232706 629778 233262 630334
rect 232706 593778 233262 594334
rect 232706 557778 233262 558334
rect 232706 521778 233262 522334
rect 232706 485778 233262 486334
rect 232706 449778 233262 450334
rect 232706 413778 233262 414334
rect 232706 377778 233262 378334
rect 232706 341778 233262 342334
rect 232706 305778 233262 306334
rect 232706 269778 233262 270334
rect 231290 255218 231526 255454
rect 231290 254898 231526 255134
rect 228986 230058 229542 230614
rect 232706 233778 233262 234334
rect 231290 219218 231526 219454
rect 231290 218898 231526 219134
rect 228986 194058 229542 194614
rect 232706 197778 233262 198334
rect 231290 183218 231526 183454
rect 231290 182898 231526 183134
rect 228986 158058 229542 158614
rect 232706 161778 233262 162334
rect 231290 147218 231526 147454
rect 231290 146898 231526 147134
rect 228986 122058 229542 122614
rect 232706 125778 233262 126334
rect 231290 111218 231526 111454
rect 231290 110898 231526 111134
rect 228986 86058 229542 86614
rect 232706 89778 233262 90334
rect 231290 75218 231526 75454
rect 231290 74898 231526 75134
rect 228986 50058 229542 50614
rect 232706 53778 233262 54334
rect 231290 39218 231526 39454
rect 231290 38898 231526 39134
rect 228986 14058 229542 14614
rect 228986 -3782 229542 -3226
rect 232706 17778 233262 18334
rect 232706 -4742 233262 -4186
rect 236426 709082 236982 709638
rect 236426 669498 236982 670054
rect 236426 633498 236982 634054
rect 236426 597498 236982 598054
rect 236426 561498 236982 562054
rect 236426 525498 236982 526054
rect 236426 489498 236982 490054
rect 236426 453498 236982 454054
rect 236426 417498 236982 418054
rect 236426 381498 236982 382054
rect 236426 345498 236982 346054
rect 236426 309498 236982 310054
rect 236426 273498 236982 274054
rect 240146 710042 240702 710598
rect 240146 673218 240702 673774
rect 240146 637218 240702 637774
rect 240146 601218 240702 601774
rect 240146 565218 240702 565774
rect 240146 529218 240702 529774
rect 240146 493218 240702 493774
rect 240146 457218 240702 457774
rect 240146 421218 240702 421774
rect 240146 385218 240702 385774
rect 240146 349218 240702 349774
rect 240146 313218 240702 313774
rect 240146 277218 240702 277774
rect 238970 258938 239206 259174
rect 238970 258618 239206 258854
rect 236426 237498 236982 238054
rect 240146 241218 240702 241774
rect 238970 222938 239206 223174
rect 238970 222618 239206 222854
rect 236426 201498 236982 202054
rect 240146 205218 240702 205774
rect 238970 186938 239206 187174
rect 238970 186618 239206 186854
rect 236426 165498 236982 166054
rect 240146 169218 240702 169774
rect 238970 150938 239206 151174
rect 238970 150618 239206 150854
rect 236426 129498 236982 130054
rect 240146 133218 240702 133774
rect 238970 114938 239206 115174
rect 238970 114618 239206 114854
rect 236426 93498 236982 94054
rect 240146 97218 240702 97774
rect 238970 78938 239206 79174
rect 238970 78618 239206 78854
rect 236426 57498 236982 58054
rect 240146 61218 240702 61774
rect 238970 42938 239206 43174
rect 238970 42618 239206 42854
rect 236426 21498 236982 22054
rect 240146 25218 240702 25774
rect 238970 6938 239206 7174
rect 238970 6618 239206 6854
rect 236426 -5702 236982 -5146
rect 240146 -6662 240702 -6106
rect 243866 711002 244422 711558
rect 243866 676938 244422 677494
rect 243866 640938 244422 641494
rect 243866 604938 244422 605494
rect 243866 568938 244422 569494
rect 243866 532938 244422 533494
rect 243866 496938 244422 497494
rect 243866 460938 244422 461494
rect 243866 424938 244422 425494
rect 243866 388938 244422 389494
rect 243866 352938 244422 353494
rect 243866 316938 244422 317494
rect 253826 704282 254382 704838
rect 253826 686898 254382 687454
rect 253826 650898 254382 651454
rect 253826 614898 254382 615454
rect 253826 578898 254382 579454
rect 253826 542898 254382 543454
rect 253826 506898 254382 507454
rect 253826 470898 254382 471454
rect 253826 434898 254382 435454
rect 253826 398898 254382 399454
rect 253826 362898 254382 363454
rect 253826 326898 254382 327454
rect 253826 290898 254382 291454
rect 257546 705242 258102 705798
rect 257546 690618 258102 691174
rect 257546 654618 258102 655174
rect 257546 618618 258102 619174
rect 257546 582618 258102 583174
rect 257546 546618 258102 547174
rect 257546 510618 258102 511174
rect 257546 474618 258102 475174
rect 257546 438618 258102 439174
rect 257546 402618 258102 403174
rect 257546 366618 258102 367174
rect 257546 330618 258102 331174
rect 257546 294618 258102 295174
rect 243866 280938 244422 281494
rect 254330 273818 254566 274054
rect 254330 273498 254566 273734
rect 246650 270098 246886 270334
rect 246650 269778 246886 270014
rect 243866 244938 244422 245494
rect 261266 706202 261822 706758
rect 261266 694338 261822 694894
rect 261266 658338 261822 658894
rect 261266 622338 261822 622894
rect 261266 586338 261822 586894
rect 261266 550338 261822 550894
rect 261266 514338 261822 514894
rect 261266 478338 261822 478894
rect 261266 442338 261822 442894
rect 261266 406338 261822 406894
rect 261266 370338 261822 370894
rect 261266 334338 261822 334894
rect 261266 298338 261822 298894
rect 264986 707162 265542 707718
rect 264986 698058 265542 698614
rect 264986 662058 265542 662614
rect 264986 626058 265542 626614
rect 264986 590058 265542 590614
rect 264986 554058 265542 554614
rect 264986 518058 265542 518614
rect 264986 482058 265542 482614
rect 264986 446058 265542 446614
rect 264986 410058 265542 410614
rect 264986 374058 265542 374614
rect 264986 338058 265542 338614
rect 264986 302058 265542 302614
rect 257546 258618 258102 259174
rect 254330 237818 254566 238054
rect 254330 237498 254566 237734
rect 246650 234098 246886 234334
rect 246650 233778 246886 234014
rect 243866 208938 244422 209494
rect 264986 266058 265542 266614
rect 262010 255218 262246 255454
rect 262010 254898 262246 255134
rect 257546 222618 258102 223174
rect 254330 201818 254566 202054
rect 254330 201498 254566 201734
rect 246650 198098 246886 198334
rect 246650 197778 246886 198014
rect 243866 172938 244422 173494
rect 264986 230058 265542 230614
rect 262010 219218 262246 219454
rect 262010 218898 262246 219134
rect 257546 186618 258102 187174
rect 254330 165818 254566 166054
rect 254330 165498 254566 165734
rect 246650 162098 246886 162334
rect 246650 161778 246886 162014
rect 243866 136938 244422 137494
rect 264986 194058 265542 194614
rect 262010 183218 262246 183454
rect 262010 182898 262246 183134
rect 257546 150618 258102 151174
rect 254330 129818 254566 130054
rect 254330 129498 254566 129734
rect 246650 126098 246886 126334
rect 246650 125778 246886 126014
rect 243866 100938 244422 101494
rect 264986 158058 265542 158614
rect 262010 147218 262246 147454
rect 262010 146898 262246 147134
rect 257546 114618 258102 115174
rect 254330 93818 254566 94054
rect 254330 93498 254566 93734
rect 246650 90098 246886 90334
rect 246650 89778 246886 90014
rect 243866 64938 244422 65494
rect 264986 122058 265542 122614
rect 262010 111218 262246 111454
rect 262010 110898 262246 111134
rect 257546 78618 258102 79174
rect 254330 57818 254566 58054
rect 254330 57498 254566 57734
rect 246650 54098 246886 54334
rect 246650 53778 246886 54014
rect 243866 28938 244422 29494
rect 264986 86058 265542 86614
rect 262010 75218 262246 75454
rect 262010 74898 262246 75134
rect 257546 42618 258102 43174
rect 254330 21818 254566 22054
rect 254330 21498 254566 21734
rect 246650 18098 246886 18334
rect 246650 17778 246886 18014
rect 264986 50058 265542 50614
rect 262010 39218 262246 39454
rect 262010 38898 262246 39134
rect 257546 6618 258102 7174
rect 243866 -7622 244422 -7066
rect 253826 -902 254382 -346
rect 264986 14058 265542 14614
rect 257546 -1862 258102 -1306
rect 261266 -2822 261822 -2266
rect 264986 -3782 265542 -3226
rect 268706 708122 269262 708678
rect 268706 665778 269262 666334
rect 268706 629778 269262 630334
rect 268706 593778 269262 594334
rect 268706 557778 269262 558334
rect 268706 521778 269262 522334
rect 268706 485778 269262 486334
rect 268706 449778 269262 450334
rect 268706 413778 269262 414334
rect 268706 377778 269262 378334
rect 268706 341778 269262 342334
rect 268706 305778 269262 306334
rect 268706 269778 269262 270334
rect 272426 709082 272982 709638
rect 272426 669498 272982 670054
rect 272426 633498 272982 634054
rect 272426 597498 272982 598054
rect 272426 561498 272982 562054
rect 272426 525498 272982 526054
rect 272426 489498 272982 490054
rect 272426 453498 272982 454054
rect 272426 417498 272982 418054
rect 272426 381498 272982 382054
rect 272426 345498 272982 346054
rect 272426 309498 272982 310054
rect 272426 273498 272982 274054
rect 269690 258938 269926 259174
rect 269690 258618 269926 258854
rect 268706 233778 269262 234334
rect 272426 237498 272982 238054
rect 269690 222938 269926 223174
rect 269690 222618 269926 222854
rect 268706 197778 269262 198334
rect 272426 201498 272982 202054
rect 269690 186938 269926 187174
rect 269690 186618 269926 186854
rect 268706 161778 269262 162334
rect 272426 165498 272982 166054
rect 269690 150938 269926 151174
rect 269690 150618 269926 150854
rect 268706 125778 269262 126334
rect 272426 129498 272982 130054
rect 269690 114938 269926 115174
rect 269690 114618 269926 114854
rect 268706 89778 269262 90334
rect 272426 93498 272982 94054
rect 269690 78938 269926 79174
rect 269690 78618 269926 78854
rect 268706 53778 269262 54334
rect 272426 57498 272982 58054
rect 269690 42938 269926 43174
rect 269690 42618 269926 42854
rect 268706 17778 269262 18334
rect 272426 21498 272982 22054
rect 269690 6938 269926 7174
rect 269690 6618 269926 6854
rect 268706 -4742 269262 -4186
rect 272426 -5702 272982 -5146
rect 276146 710042 276702 710598
rect 276146 673218 276702 673774
rect 276146 637218 276702 637774
rect 276146 601218 276702 601774
rect 276146 565218 276702 565774
rect 276146 529218 276702 529774
rect 276146 493218 276702 493774
rect 276146 457218 276702 457774
rect 276146 421218 276702 421774
rect 276146 385218 276702 385774
rect 276146 349218 276702 349774
rect 276146 313218 276702 313774
rect 276146 277218 276702 277774
rect 279866 711002 280422 711558
rect 279866 676938 280422 677494
rect 279866 640938 280422 641494
rect 279866 604938 280422 605494
rect 279866 568938 280422 569494
rect 279866 532938 280422 533494
rect 279866 496938 280422 497494
rect 279866 460938 280422 461494
rect 279866 424938 280422 425494
rect 279866 388938 280422 389494
rect 279866 352938 280422 353494
rect 279866 316938 280422 317494
rect 279866 280938 280422 281494
rect 277370 270098 277606 270334
rect 277370 269778 277606 270014
rect 276146 241218 276702 241774
rect 289826 704282 290382 704838
rect 289826 686898 290382 687454
rect 289826 650898 290382 651454
rect 289826 614898 290382 615454
rect 289826 578898 290382 579454
rect 289826 542898 290382 543454
rect 289826 506898 290382 507454
rect 289826 470898 290382 471454
rect 289826 434898 290382 435454
rect 289826 398898 290382 399454
rect 289826 362898 290382 363454
rect 289826 326898 290382 327454
rect 289826 290898 290382 291454
rect 285050 273818 285286 274054
rect 285050 273498 285286 273734
rect 279866 244938 280422 245494
rect 277370 234098 277606 234334
rect 277370 233778 277606 234014
rect 276146 205218 276702 205774
rect 289826 254898 290382 255454
rect 285050 237818 285286 238054
rect 285050 237498 285286 237734
rect 279866 208938 280422 209494
rect 277370 198098 277606 198334
rect 277370 197778 277606 198014
rect 276146 169218 276702 169774
rect 289826 218898 290382 219454
rect 285050 201818 285286 202054
rect 285050 201498 285286 201734
rect 279866 172938 280422 173494
rect 277370 162098 277606 162334
rect 277370 161778 277606 162014
rect 276146 133218 276702 133774
rect 289826 182898 290382 183454
rect 285050 165818 285286 166054
rect 285050 165498 285286 165734
rect 279866 136938 280422 137494
rect 277370 126098 277606 126334
rect 277370 125778 277606 126014
rect 276146 97218 276702 97774
rect 289826 146898 290382 147454
rect 285050 129818 285286 130054
rect 285050 129498 285286 129734
rect 279866 100938 280422 101494
rect 277370 90098 277606 90334
rect 277370 89778 277606 90014
rect 276146 61218 276702 61774
rect 289826 110898 290382 111454
rect 285050 93818 285286 94054
rect 285050 93498 285286 93734
rect 279866 64938 280422 65494
rect 277370 54098 277606 54334
rect 277370 53778 277606 54014
rect 276146 25218 276702 25774
rect 289826 74898 290382 75454
rect 285050 57818 285286 58054
rect 285050 57498 285286 57734
rect 279866 28938 280422 29494
rect 277370 18098 277606 18334
rect 277370 17778 277606 18014
rect 276146 -6662 276702 -6106
rect 289826 38898 290382 39454
rect 285050 21818 285286 22054
rect 285050 21498 285286 21734
rect 279866 -7622 280422 -7066
rect 289826 2898 290382 3454
rect 289826 -902 290382 -346
rect 293546 705242 294102 705798
rect 293546 690618 294102 691174
rect 293546 654618 294102 655174
rect 293546 618618 294102 619174
rect 293546 582618 294102 583174
rect 293546 546618 294102 547174
rect 293546 510618 294102 511174
rect 293546 474618 294102 475174
rect 293546 438618 294102 439174
rect 293546 402618 294102 403174
rect 293546 366618 294102 367174
rect 293546 330618 294102 331174
rect 293546 294618 294102 295174
rect 293546 258618 294102 259174
rect 293546 222618 294102 223174
rect 293546 186618 294102 187174
rect 293546 150618 294102 151174
rect 293546 114618 294102 115174
rect 293546 78618 294102 79174
rect 293546 42618 294102 43174
rect 293546 6618 294102 7174
rect 293546 -1862 294102 -1306
rect 297266 706202 297822 706758
rect 297266 694338 297822 694894
rect 297266 658338 297822 658894
rect 297266 622338 297822 622894
rect 297266 586338 297822 586894
rect 297266 550338 297822 550894
rect 297266 514338 297822 514894
rect 297266 478338 297822 478894
rect 297266 442338 297822 442894
rect 297266 406338 297822 406894
rect 297266 370338 297822 370894
rect 297266 334338 297822 334894
rect 297266 298338 297822 298894
rect 297266 262338 297822 262894
rect 297266 226338 297822 226894
rect 297266 190338 297822 190894
rect 297266 154338 297822 154894
rect 297266 118338 297822 118894
rect 297266 82338 297822 82894
rect 297266 46338 297822 46894
rect 297266 10338 297822 10894
rect 297266 -2822 297822 -2266
rect 300986 707162 301542 707718
rect 300986 698058 301542 698614
rect 300986 662058 301542 662614
rect 300986 626058 301542 626614
rect 300986 590058 301542 590614
rect 300986 554058 301542 554614
rect 300986 518058 301542 518614
rect 300986 482058 301542 482614
rect 300986 446058 301542 446614
rect 300986 410058 301542 410614
rect 300986 374058 301542 374614
rect 300986 338058 301542 338614
rect 300986 302058 301542 302614
rect 300986 266058 301542 266614
rect 300986 230058 301542 230614
rect 300986 194058 301542 194614
rect 300986 158058 301542 158614
rect 300986 122058 301542 122614
rect 300986 86058 301542 86614
rect 300986 50058 301542 50614
rect 300986 14058 301542 14614
rect 300986 -3782 301542 -3226
rect 304706 708122 305262 708678
rect 304706 665778 305262 666334
rect 304706 629778 305262 630334
rect 304706 593778 305262 594334
rect 304706 557778 305262 558334
rect 304706 521778 305262 522334
rect 304706 485778 305262 486334
rect 304706 449778 305262 450334
rect 304706 413778 305262 414334
rect 304706 377778 305262 378334
rect 304706 341778 305262 342334
rect 304706 305778 305262 306334
rect 304706 269778 305262 270334
rect 304706 233778 305262 234334
rect 304706 197778 305262 198334
rect 304706 161778 305262 162334
rect 304706 125778 305262 126334
rect 304706 89778 305262 90334
rect 304706 53778 305262 54334
rect 304706 17778 305262 18334
rect 304706 -4742 305262 -4186
rect 308426 709082 308982 709638
rect 308426 669498 308982 670054
rect 308426 633498 308982 634054
rect 308426 597498 308982 598054
rect 308426 561498 308982 562054
rect 308426 525498 308982 526054
rect 308426 489498 308982 490054
rect 308426 453498 308982 454054
rect 308426 417498 308982 418054
rect 308426 381498 308982 382054
rect 308426 345498 308982 346054
rect 308426 309498 308982 310054
rect 308426 273498 308982 274054
rect 308426 237498 308982 238054
rect 308426 201498 308982 202054
rect 308426 165498 308982 166054
rect 308426 129498 308982 130054
rect 308426 93498 308982 94054
rect 308426 57498 308982 58054
rect 308426 21498 308982 22054
rect 308426 -5702 308982 -5146
rect 312146 710042 312702 710598
rect 312146 673218 312702 673774
rect 312146 637218 312702 637774
rect 312146 601218 312702 601774
rect 312146 565218 312702 565774
rect 312146 529218 312702 529774
rect 312146 493218 312702 493774
rect 312146 457218 312702 457774
rect 312146 421218 312702 421774
rect 312146 385218 312702 385774
rect 312146 349218 312702 349774
rect 312146 313218 312702 313774
rect 312146 277218 312702 277774
rect 312146 241218 312702 241774
rect 312146 205218 312702 205774
rect 312146 169218 312702 169774
rect 312146 133218 312702 133774
rect 312146 97218 312702 97774
rect 312146 61218 312702 61774
rect 312146 25218 312702 25774
rect 312146 -6662 312702 -6106
rect 315866 711002 316422 711558
rect 315866 676938 316422 677494
rect 315866 640938 316422 641494
rect 315866 604938 316422 605494
rect 315866 568938 316422 569494
rect 315866 532938 316422 533494
rect 315866 496938 316422 497494
rect 315866 460938 316422 461494
rect 315866 424938 316422 425494
rect 315866 388938 316422 389494
rect 315866 352938 316422 353494
rect 315866 316938 316422 317494
rect 315866 280938 316422 281494
rect 315866 244938 316422 245494
rect 315866 208938 316422 209494
rect 315866 172938 316422 173494
rect 315866 136938 316422 137494
rect 315866 100938 316422 101494
rect 315866 64938 316422 65494
rect 315866 28938 316422 29494
rect 315866 -7622 316422 -7066
rect 325826 704282 326382 704838
rect 325826 686898 326382 687454
rect 325826 650898 326382 651454
rect 325826 614898 326382 615454
rect 325826 578898 326382 579454
rect 325826 542898 326382 543454
rect 325826 506898 326382 507454
rect 325826 470898 326382 471454
rect 325826 434898 326382 435454
rect 325826 398898 326382 399454
rect 325826 362898 326382 363454
rect 325826 326898 326382 327454
rect 325826 290898 326382 291454
rect 325826 254898 326382 255454
rect 325826 218898 326382 219454
rect 325826 182898 326382 183454
rect 325826 146898 326382 147454
rect 325826 110898 326382 111454
rect 325826 74898 326382 75454
rect 325826 38898 326382 39454
rect 325826 2898 326382 3454
rect 325826 -902 326382 -346
rect 329546 705242 330102 705798
rect 329546 690618 330102 691174
rect 329546 654618 330102 655174
rect 329546 618618 330102 619174
rect 329546 582618 330102 583174
rect 329546 546618 330102 547174
rect 329546 510618 330102 511174
rect 329546 474618 330102 475174
rect 329546 438618 330102 439174
rect 329546 402618 330102 403174
rect 329546 366618 330102 367174
rect 329546 330618 330102 331174
rect 329546 294618 330102 295174
rect 329546 258618 330102 259174
rect 329546 222618 330102 223174
rect 329546 186618 330102 187174
rect 329546 150618 330102 151174
rect 329546 114618 330102 115174
rect 329546 78618 330102 79174
rect 329546 42618 330102 43174
rect 329546 6618 330102 7174
rect 329546 -1862 330102 -1306
rect 333266 706202 333822 706758
rect 333266 694338 333822 694894
rect 333266 658338 333822 658894
rect 333266 622338 333822 622894
rect 333266 586338 333822 586894
rect 333266 550338 333822 550894
rect 333266 514338 333822 514894
rect 333266 478338 333822 478894
rect 333266 442338 333822 442894
rect 333266 406338 333822 406894
rect 333266 370338 333822 370894
rect 333266 334338 333822 334894
rect 333266 298338 333822 298894
rect 333266 262338 333822 262894
rect 333266 226338 333822 226894
rect 333266 190338 333822 190894
rect 333266 154338 333822 154894
rect 333266 118338 333822 118894
rect 333266 82338 333822 82894
rect 333266 46338 333822 46894
rect 333266 10338 333822 10894
rect 333266 -2822 333822 -2266
rect 336986 707162 337542 707718
rect 336986 698058 337542 698614
rect 336986 662058 337542 662614
rect 336986 626058 337542 626614
rect 336986 590058 337542 590614
rect 336986 554058 337542 554614
rect 336986 518058 337542 518614
rect 336986 482058 337542 482614
rect 336986 446058 337542 446614
rect 336986 410058 337542 410614
rect 336986 374058 337542 374614
rect 336986 338058 337542 338614
rect 336986 302058 337542 302614
rect 336986 266058 337542 266614
rect 336986 230058 337542 230614
rect 336986 194058 337542 194614
rect 336986 158058 337542 158614
rect 336986 122058 337542 122614
rect 336986 86058 337542 86614
rect 336986 50058 337542 50614
rect 336986 14058 337542 14614
rect 336986 -3782 337542 -3226
rect 340706 708122 341262 708678
rect 340706 665778 341262 666334
rect 340706 629778 341262 630334
rect 340706 593778 341262 594334
rect 340706 557778 341262 558334
rect 340706 521778 341262 522334
rect 340706 485778 341262 486334
rect 340706 449778 341262 450334
rect 340706 413778 341262 414334
rect 340706 377778 341262 378334
rect 340706 341778 341262 342334
rect 340706 305778 341262 306334
rect 340706 269778 341262 270334
rect 340706 233778 341262 234334
rect 340706 197778 341262 198334
rect 340706 161778 341262 162334
rect 340706 125778 341262 126334
rect 340706 89778 341262 90334
rect 340706 53778 341262 54334
rect 340706 17778 341262 18334
rect 340706 -4742 341262 -4186
rect 344426 709082 344982 709638
rect 344426 669498 344982 670054
rect 344426 633498 344982 634054
rect 344426 597498 344982 598054
rect 344426 561498 344982 562054
rect 344426 525498 344982 526054
rect 344426 489498 344982 490054
rect 344426 453498 344982 454054
rect 344426 417498 344982 418054
rect 344426 381498 344982 382054
rect 344426 345498 344982 346054
rect 344426 309498 344982 310054
rect 344426 273498 344982 274054
rect 344426 237498 344982 238054
rect 344426 201498 344982 202054
rect 344426 165498 344982 166054
rect 344426 129498 344982 130054
rect 344426 93498 344982 94054
rect 344426 57498 344982 58054
rect 344426 21498 344982 22054
rect 344426 -5702 344982 -5146
rect 348146 710042 348702 710598
rect 348146 673218 348702 673774
rect 348146 637218 348702 637774
rect 348146 601218 348702 601774
rect 348146 565218 348702 565774
rect 348146 529218 348702 529774
rect 348146 493218 348702 493774
rect 348146 457218 348702 457774
rect 348146 421218 348702 421774
rect 348146 385218 348702 385774
rect 348146 349218 348702 349774
rect 348146 313218 348702 313774
rect 348146 277218 348702 277774
rect 348146 241218 348702 241774
rect 348146 205218 348702 205774
rect 348146 169218 348702 169774
rect 348146 133218 348702 133774
rect 348146 97218 348702 97774
rect 348146 61218 348702 61774
rect 348146 25218 348702 25774
rect 348146 -6662 348702 -6106
rect 351866 711002 352422 711558
rect 351866 676938 352422 677494
rect 351866 640938 352422 641494
rect 351866 604938 352422 605494
rect 351866 568938 352422 569494
rect 351866 532938 352422 533494
rect 351866 496938 352422 497494
rect 351866 460938 352422 461494
rect 351866 424938 352422 425494
rect 351866 388938 352422 389494
rect 351866 352938 352422 353494
rect 351866 316938 352422 317494
rect 351866 280938 352422 281494
rect 351866 244938 352422 245494
rect 351866 208938 352422 209494
rect 351866 172938 352422 173494
rect 351866 136938 352422 137494
rect 351866 100938 352422 101494
rect 351866 64938 352422 65494
rect 351866 28938 352422 29494
rect 351866 -7622 352422 -7066
rect 361826 704282 362382 704838
rect 361826 686898 362382 687454
rect 361826 650898 362382 651454
rect 361826 614898 362382 615454
rect 361826 578898 362382 579454
rect 361826 542898 362382 543454
rect 361826 506898 362382 507454
rect 361826 470898 362382 471454
rect 361826 434898 362382 435454
rect 361826 398898 362382 399454
rect 361826 362898 362382 363454
rect 361826 326898 362382 327454
rect 361826 290898 362382 291454
rect 361826 254898 362382 255454
rect 361826 218898 362382 219454
rect 361826 182898 362382 183454
rect 361826 146898 362382 147454
rect 361826 110898 362382 111454
rect 361826 74898 362382 75454
rect 361826 38898 362382 39454
rect 361826 2898 362382 3454
rect 361826 -902 362382 -346
rect 365546 705242 366102 705798
rect 365546 690618 366102 691174
rect 365546 654618 366102 655174
rect 365546 618618 366102 619174
rect 365546 582618 366102 583174
rect 365546 546618 366102 547174
rect 365546 510618 366102 511174
rect 365546 474618 366102 475174
rect 365546 438618 366102 439174
rect 365546 402618 366102 403174
rect 365546 366618 366102 367174
rect 365546 330618 366102 331174
rect 365546 294618 366102 295174
rect 365546 258618 366102 259174
rect 365546 222618 366102 223174
rect 365546 186618 366102 187174
rect 365546 150618 366102 151174
rect 365546 114618 366102 115174
rect 365546 78618 366102 79174
rect 365546 42618 366102 43174
rect 365546 6618 366102 7174
rect 365546 -1862 366102 -1306
rect 369266 706202 369822 706758
rect 369266 694338 369822 694894
rect 369266 658338 369822 658894
rect 369266 622338 369822 622894
rect 369266 586338 369822 586894
rect 369266 550338 369822 550894
rect 369266 514338 369822 514894
rect 369266 478338 369822 478894
rect 369266 442338 369822 442894
rect 369266 406338 369822 406894
rect 369266 370338 369822 370894
rect 369266 334338 369822 334894
rect 369266 298338 369822 298894
rect 369266 262338 369822 262894
rect 369266 226338 369822 226894
rect 369266 190338 369822 190894
rect 369266 154338 369822 154894
rect 369266 118338 369822 118894
rect 369266 82338 369822 82894
rect 369266 46338 369822 46894
rect 369266 10338 369822 10894
rect 369266 -2822 369822 -2266
rect 372986 707162 373542 707718
rect 372986 698058 373542 698614
rect 372986 662058 373542 662614
rect 372986 626058 373542 626614
rect 372986 590058 373542 590614
rect 372986 554058 373542 554614
rect 372986 518058 373542 518614
rect 372986 482058 373542 482614
rect 372986 446058 373542 446614
rect 372986 410058 373542 410614
rect 372986 374058 373542 374614
rect 372986 338058 373542 338614
rect 372986 302058 373542 302614
rect 372986 266058 373542 266614
rect 372986 230058 373542 230614
rect 372986 194058 373542 194614
rect 372986 158058 373542 158614
rect 372986 122058 373542 122614
rect 372986 86058 373542 86614
rect 372986 50058 373542 50614
rect 372986 14058 373542 14614
rect 372986 -3782 373542 -3226
rect 376706 708122 377262 708678
rect 376706 665778 377262 666334
rect 376706 629778 377262 630334
rect 376706 593778 377262 594334
rect 376706 557778 377262 558334
rect 376706 521778 377262 522334
rect 376706 485778 377262 486334
rect 376706 449778 377262 450334
rect 376706 413778 377262 414334
rect 376706 377778 377262 378334
rect 376706 341778 377262 342334
rect 376706 305778 377262 306334
rect 376706 269778 377262 270334
rect 376706 233778 377262 234334
rect 376706 197778 377262 198334
rect 376706 161778 377262 162334
rect 376706 125778 377262 126334
rect 376706 89778 377262 90334
rect 376706 53778 377262 54334
rect 376706 17778 377262 18334
rect 376706 -4742 377262 -4186
rect 380426 709082 380982 709638
rect 380426 669498 380982 670054
rect 380426 633498 380982 634054
rect 380426 597498 380982 598054
rect 380426 561498 380982 562054
rect 380426 525498 380982 526054
rect 380426 489498 380982 490054
rect 380426 453498 380982 454054
rect 380426 417498 380982 418054
rect 380426 381498 380982 382054
rect 380426 345498 380982 346054
rect 380426 309498 380982 310054
rect 380426 273498 380982 274054
rect 380426 237498 380982 238054
rect 380426 201498 380982 202054
rect 380426 165498 380982 166054
rect 380426 129498 380982 130054
rect 380426 93498 380982 94054
rect 380426 57498 380982 58054
rect 380426 21498 380982 22054
rect 380426 -5702 380982 -5146
rect 384146 710042 384702 710598
rect 384146 673218 384702 673774
rect 384146 637218 384702 637774
rect 384146 601218 384702 601774
rect 384146 565218 384702 565774
rect 384146 529218 384702 529774
rect 384146 493218 384702 493774
rect 384146 457218 384702 457774
rect 384146 421218 384702 421774
rect 384146 385218 384702 385774
rect 384146 349218 384702 349774
rect 384146 313218 384702 313774
rect 384146 277218 384702 277774
rect 384146 241218 384702 241774
rect 384146 205218 384702 205774
rect 384146 169218 384702 169774
rect 384146 133218 384702 133774
rect 384146 97218 384702 97774
rect 384146 61218 384702 61774
rect 384146 25218 384702 25774
rect 384146 -6662 384702 -6106
rect 387866 711002 388422 711558
rect 387866 676938 388422 677494
rect 387866 640938 388422 641494
rect 387866 604938 388422 605494
rect 387866 568938 388422 569494
rect 387866 532938 388422 533494
rect 387866 496938 388422 497494
rect 387866 460938 388422 461494
rect 387866 424938 388422 425494
rect 387866 388938 388422 389494
rect 387866 352938 388422 353494
rect 387866 316938 388422 317494
rect 387866 280938 388422 281494
rect 387866 244938 388422 245494
rect 387866 208938 388422 209494
rect 387866 172938 388422 173494
rect 387866 136938 388422 137494
rect 387866 100938 388422 101494
rect 387866 64938 388422 65494
rect 387866 28938 388422 29494
rect 387866 -7622 388422 -7066
rect 397826 704282 398382 704838
rect 397826 686898 398382 687454
rect 397826 650898 398382 651454
rect 397826 614898 398382 615454
rect 397826 578898 398382 579454
rect 397826 542898 398382 543454
rect 397826 506898 398382 507454
rect 397826 470898 398382 471454
rect 397826 434898 398382 435454
rect 397826 398898 398382 399454
rect 397826 362898 398382 363454
rect 397826 326898 398382 327454
rect 397826 290898 398382 291454
rect 397826 254898 398382 255454
rect 397826 218898 398382 219454
rect 397826 182898 398382 183454
rect 397826 146898 398382 147454
rect 397826 110898 398382 111454
rect 397826 74898 398382 75454
rect 397826 38898 398382 39454
rect 397826 2898 398382 3454
rect 397826 -902 398382 -346
rect 401546 705242 402102 705798
rect 401546 690618 402102 691174
rect 401546 654618 402102 655174
rect 401546 618618 402102 619174
rect 401546 582618 402102 583174
rect 401546 546618 402102 547174
rect 401546 510618 402102 511174
rect 401546 474618 402102 475174
rect 401546 438618 402102 439174
rect 401546 402618 402102 403174
rect 401546 366618 402102 367174
rect 401546 330618 402102 331174
rect 401546 294618 402102 295174
rect 401546 258618 402102 259174
rect 401546 222618 402102 223174
rect 401546 186618 402102 187174
rect 401546 150618 402102 151174
rect 401546 114618 402102 115174
rect 401546 78618 402102 79174
rect 401546 42618 402102 43174
rect 401546 6618 402102 7174
rect 401546 -1862 402102 -1306
rect 405266 706202 405822 706758
rect 405266 694338 405822 694894
rect 405266 658338 405822 658894
rect 405266 622338 405822 622894
rect 405266 586338 405822 586894
rect 405266 550338 405822 550894
rect 405266 514338 405822 514894
rect 405266 478338 405822 478894
rect 405266 442338 405822 442894
rect 405266 406338 405822 406894
rect 405266 370338 405822 370894
rect 405266 334338 405822 334894
rect 405266 298338 405822 298894
rect 405266 262338 405822 262894
rect 405266 226338 405822 226894
rect 405266 190338 405822 190894
rect 405266 154338 405822 154894
rect 405266 118338 405822 118894
rect 405266 82338 405822 82894
rect 405266 46338 405822 46894
rect 405266 10338 405822 10894
rect 405266 -2822 405822 -2266
rect 408986 707162 409542 707718
rect 408986 698058 409542 698614
rect 408986 662058 409542 662614
rect 408986 626058 409542 626614
rect 408986 590058 409542 590614
rect 408986 554058 409542 554614
rect 408986 518058 409542 518614
rect 408986 482058 409542 482614
rect 408986 446058 409542 446614
rect 408986 410058 409542 410614
rect 408986 374058 409542 374614
rect 408986 338058 409542 338614
rect 408986 302058 409542 302614
rect 408986 266058 409542 266614
rect 408986 230058 409542 230614
rect 408986 194058 409542 194614
rect 408986 158058 409542 158614
rect 408986 122058 409542 122614
rect 408986 86058 409542 86614
rect 408986 50058 409542 50614
rect 408986 14058 409542 14614
rect 408986 -3782 409542 -3226
rect 412706 708122 413262 708678
rect 412706 665778 413262 666334
rect 412706 629778 413262 630334
rect 412706 593778 413262 594334
rect 412706 557778 413262 558334
rect 412706 521778 413262 522334
rect 412706 485778 413262 486334
rect 412706 449778 413262 450334
rect 412706 413778 413262 414334
rect 412706 377778 413262 378334
rect 412706 341778 413262 342334
rect 412706 305778 413262 306334
rect 412706 269778 413262 270334
rect 412706 233778 413262 234334
rect 412706 197778 413262 198334
rect 412706 161778 413262 162334
rect 412706 125778 413262 126334
rect 412706 89778 413262 90334
rect 412706 53778 413262 54334
rect 412706 17778 413262 18334
rect 412706 -4742 413262 -4186
rect 416426 709082 416982 709638
rect 416426 669498 416982 670054
rect 416426 633498 416982 634054
rect 416426 597498 416982 598054
rect 416426 561498 416982 562054
rect 416426 525498 416982 526054
rect 416426 489498 416982 490054
rect 416426 453498 416982 454054
rect 416426 417498 416982 418054
rect 416426 381498 416982 382054
rect 416426 345498 416982 346054
rect 416426 309498 416982 310054
rect 416426 273498 416982 274054
rect 416426 237498 416982 238054
rect 416426 201498 416982 202054
rect 416426 165498 416982 166054
rect 416426 129498 416982 130054
rect 416426 93498 416982 94054
rect 416426 57498 416982 58054
rect 416426 21498 416982 22054
rect 416426 -5702 416982 -5146
rect 420146 710042 420702 710598
rect 420146 673218 420702 673774
rect 420146 637218 420702 637774
rect 420146 601218 420702 601774
rect 420146 565218 420702 565774
rect 420146 529218 420702 529774
rect 420146 493218 420702 493774
rect 420146 457218 420702 457774
rect 420146 421218 420702 421774
rect 420146 385218 420702 385774
rect 420146 349218 420702 349774
rect 420146 313218 420702 313774
rect 420146 277218 420702 277774
rect 420146 241218 420702 241774
rect 420146 205218 420702 205774
rect 420146 169218 420702 169774
rect 420146 133218 420702 133774
rect 420146 97218 420702 97774
rect 420146 61218 420702 61774
rect 420146 25218 420702 25774
rect 420146 -6662 420702 -6106
rect 423866 711002 424422 711558
rect 423866 676938 424422 677494
rect 423866 640938 424422 641494
rect 423866 604938 424422 605494
rect 423866 568938 424422 569494
rect 423866 532938 424422 533494
rect 423866 496938 424422 497494
rect 423866 460938 424422 461494
rect 423866 424938 424422 425494
rect 423866 388938 424422 389494
rect 423866 352938 424422 353494
rect 423866 316938 424422 317494
rect 423866 280938 424422 281494
rect 423866 244938 424422 245494
rect 423866 208938 424422 209494
rect 423866 172938 424422 173494
rect 423866 136938 424422 137494
rect 423866 100938 424422 101494
rect 423866 64938 424422 65494
rect 423866 28938 424422 29494
rect 423866 -7622 424422 -7066
rect 433826 704282 434382 704838
rect 433826 686898 434382 687454
rect 433826 650898 434382 651454
rect 433826 614898 434382 615454
rect 433826 578898 434382 579454
rect 433826 542898 434382 543454
rect 433826 506898 434382 507454
rect 433826 470898 434382 471454
rect 433826 434898 434382 435454
rect 433826 398898 434382 399454
rect 433826 362898 434382 363454
rect 433826 326898 434382 327454
rect 433826 290898 434382 291454
rect 433826 254898 434382 255454
rect 433826 218898 434382 219454
rect 433826 182898 434382 183454
rect 433826 146898 434382 147454
rect 433826 110898 434382 111454
rect 433826 74898 434382 75454
rect 433826 38898 434382 39454
rect 433826 2898 434382 3454
rect 433826 -902 434382 -346
rect 437546 705242 438102 705798
rect 437546 690618 438102 691174
rect 437546 654618 438102 655174
rect 437546 618618 438102 619174
rect 437546 582618 438102 583174
rect 437546 546618 438102 547174
rect 437546 510618 438102 511174
rect 437546 474618 438102 475174
rect 437546 438618 438102 439174
rect 437546 402618 438102 403174
rect 437546 366618 438102 367174
rect 437546 330618 438102 331174
rect 437546 294618 438102 295174
rect 437546 258618 438102 259174
rect 437546 222618 438102 223174
rect 437546 186618 438102 187174
rect 437546 150618 438102 151174
rect 437546 114618 438102 115174
rect 437546 78618 438102 79174
rect 437546 42618 438102 43174
rect 437546 6618 438102 7174
rect 437546 -1862 438102 -1306
rect 441266 706202 441822 706758
rect 441266 694338 441822 694894
rect 441266 658338 441822 658894
rect 441266 622338 441822 622894
rect 441266 586338 441822 586894
rect 441266 550338 441822 550894
rect 441266 514338 441822 514894
rect 441266 478338 441822 478894
rect 441266 442338 441822 442894
rect 441266 406338 441822 406894
rect 441266 370338 441822 370894
rect 441266 334338 441822 334894
rect 441266 298338 441822 298894
rect 441266 262338 441822 262894
rect 441266 226338 441822 226894
rect 441266 190338 441822 190894
rect 441266 154338 441822 154894
rect 441266 118338 441822 118894
rect 441266 82338 441822 82894
rect 441266 46338 441822 46894
rect 441266 10338 441822 10894
rect 441266 -2822 441822 -2266
rect 444986 707162 445542 707718
rect 444986 698058 445542 698614
rect 444986 662058 445542 662614
rect 444986 626058 445542 626614
rect 444986 590058 445542 590614
rect 444986 554058 445542 554614
rect 444986 518058 445542 518614
rect 444986 482058 445542 482614
rect 444986 446058 445542 446614
rect 444986 410058 445542 410614
rect 444986 374058 445542 374614
rect 444986 338058 445542 338614
rect 444986 302058 445542 302614
rect 444986 266058 445542 266614
rect 444986 230058 445542 230614
rect 444986 194058 445542 194614
rect 444986 158058 445542 158614
rect 444986 122058 445542 122614
rect 444986 86058 445542 86614
rect 444986 50058 445542 50614
rect 444986 14058 445542 14614
rect 444986 -3782 445542 -3226
rect 448706 708122 449262 708678
rect 448706 665778 449262 666334
rect 448706 629778 449262 630334
rect 448706 593778 449262 594334
rect 448706 557778 449262 558334
rect 448706 521778 449262 522334
rect 448706 485778 449262 486334
rect 448706 449778 449262 450334
rect 448706 413778 449262 414334
rect 448706 377778 449262 378334
rect 448706 341778 449262 342334
rect 448706 305778 449262 306334
rect 448706 269778 449262 270334
rect 448706 233778 449262 234334
rect 448706 197778 449262 198334
rect 448706 161778 449262 162334
rect 448706 125778 449262 126334
rect 448706 89778 449262 90334
rect 448706 53778 449262 54334
rect 448706 17778 449262 18334
rect 448706 -4742 449262 -4186
rect 452426 709082 452982 709638
rect 452426 669498 452982 670054
rect 452426 633498 452982 634054
rect 452426 597498 452982 598054
rect 452426 561498 452982 562054
rect 452426 525498 452982 526054
rect 452426 489498 452982 490054
rect 452426 453498 452982 454054
rect 452426 417498 452982 418054
rect 452426 381498 452982 382054
rect 452426 345498 452982 346054
rect 452426 309498 452982 310054
rect 452426 273498 452982 274054
rect 452426 237498 452982 238054
rect 452426 201498 452982 202054
rect 452426 165498 452982 166054
rect 452426 129498 452982 130054
rect 452426 93498 452982 94054
rect 452426 57498 452982 58054
rect 452426 21498 452982 22054
rect 452426 -5702 452982 -5146
rect 456146 710042 456702 710598
rect 456146 673218 456702 673774
rect 456146 637218 456702 637774
rect 456146 601218 456702 601774
rect 456146 565218 456702 565774
rect 456146 529218 456702 529774
rect 456146 493218 456702 493774
rect 456146 457218 456702 457774
rect 456146 421218 456702 421774
rect 456146 385218 456702 385774
rect 456146 349218 456702 349774
rect 456146 313218 456702 313774
rect 456146 277218 456702 277774
rect 456146 241218 456702 241774
rect 456146 205218 456702 205774
rect 456146 169218 456702 169774
rect 456146 133218 456702 133774
rect 456146 97218 456702 97774
rect 456146 61218 456702 61774
rect 456146 25218 456702 25774
rect 456146 -6662 456702 -6106
rect 459866 711002 460422 711558
rect 459866 676938 460422 677494
rect 459866 640938 460422 641494
rect 459866 604938 460422 605494
rect 459866 568938 460422 569494
rect 459866 532938 460422 533494
rect 459866 496938 460422 497494
rect 459866 460938 460422 461494
rect 459866 424938 460422 425494
rect 459866 388938 460422 389494
rect 459866 352938 460422 353494
rect 459866 316938 460422 317494
rect 459866 280938 460422 281494
rect 459866 244938 460422 245494
rect 459866 208938 460422 209494
rect 459866 172938 460422 173494
rect 459866 136938 460422 137494
rect 459866 100938 460422 101494
rect 459866 64938 460422 65494
rect 459866 28938 460422 29494
rect 459866 -7622 460422 -7066
rect 469826 704282 470382 704838
rect 469826 686898 470382 687454
rect 469826 650898 470382 651454
rect 469826 614898 470382 615454
rect 469826 578898 470382 579454
rect 469826 542898 470382 543454
rect 469826 506898 470382 507454
rect 469826 470898 470382 471454
rect 469826 434898 470382 435454
rect 469826 398898 470382 399454
rect 469826 362898 470382 363454
rect 469826 326898 470382 327454
rect 469826 290898 470382 291454
rect 469826 254898 470382 255454
rect 469826 218898 470382 219454
rect 469826 182898 470382 183454
rect 469826 146898 470382 147454
rect 469826 110898 470382 111454
rect 469826 74898 470382 75454
rect 469826 38898 470382 39454
rect 469826 2898 470382 3454
rect 469826 -902 470382 -346
rect 473546 705242 474102 705798
rect 473546 690618 474102 691174
rect 473546 654618 474102 655174
rect 473546 618618 474102 619174
rect 473546 582618 474102 583174
rect 473546 546618 474102 547174
rect 473546 510618 474102 511174
rect 473546 474618 474102 475174
rect 473546 438618 474102 439174
rect 473546 402618 474102 403174
rect 473546 366618 474102 367174
rect 473546 330618 474102 331174
rect 473546 294618 474102 295174
rect 473546 258618 474102 259174
rect 473546 222618 474102 223174
rect 473546 186618 474102 187174
rect 473546 150618 474102 151174
rect 473546 114618 474102 115174
rect 473546 78618 474102 79174
rect 473546 42618 474102 43174
rect 473546 6618 474102 7174
rect 473546 -1862 474102 -1306
rect 477266 706202 477822 706758
rect 477266 694338 477822 694894
rect 477266 658338 477822 658894
rect 477266 622338 477822 622894
rect 477266 586338 477822 586894
rect 477266 550338 477822 550894
rect 477266 514338 477822 514894
rect 477266 478338 477822 478894
rect 477266 442338 477822 442894
rect 477266 406338 477822 406894
rect 477266 370338 477822 370894
rect 477266 334338 477822 334894
rect 477266 298338 477822 298894
rect 477266 262338 477822 262894
rect 477266 226338 477822 226894
rect 477266 190338 477822 190894
rect 477266 154338 477822 154894
rect 477266 118338 477822 118894
rect 477266 82338 477822 82894
rect 477266 46338 477822 46894
rect 477266 10338 477822 10894
rect 477266 -2822 477822 -2266
rect 480986 707162 481542 707718
rect 480986 698058 481542 698614
rect 480986 662058 481542 662614
rect 480986 626058 481542 626614
rect 480986 590058 481542 590614
rect 480986 554058 481542 554614
rect 480986 518058 481542 518614
rect 480986 482058 481542 482614
rect 480986 446058 481542 446614
rect 480986 410058 481542 410614
rect 480986 374058 481542 374614
rect 480986 338058 481542 338614
rect 480986 302058 481542 302614
rect 480986 266058 481542 266614
rect 480986 230058 481542 230614
rect 480986 194058 481542 194614
rect 480986 158058 481542 158614
rect 480986 122058 481542 122614
rect 480986 86058 481542 86614
rect 480986 50058 481542 50614
rect 480986 14058 481542 14614
rect 480986 -3782 481542 -3226
rect 484706 708122 485262 708678
rect 484706 665778 485262 666334
rect 484706 629778 485262 630334
rect 484706 593778 485262 594334
rect 484706 557778 485262 558334
rect 484706 521778 485262 522334
rect 484706 485778 485262 486334
rect 484706 449778 485262 450334
rect 484706 413778 485262 414334
rect 484706 377778 485262 378334
rect 484706 341778 485262 342334
rect 484706 305778 485262 306334
rect 484706 269778 485262 270334
rect 484706 233778 485262 234334
rect 484706 197778 485262 198334
rect 484706 161778 485262 162334
rect 484706 125778 485262 126334
rect 484706 89778 485262 90334
rect 484706 53778 485262 54334
rect 484706 17778 485262 18334
rect 484706 -4742 485262 -4186
rect 488426 709082 488982 709638
rect 488426 669498 488982 670054
rect 488426 633498 488982 634054
rect 488426 597498 488982 598054
rect 488426 561498 488982 562054
rect 488426 525498 488982 526054
rect 488426 489498 488982 490054
rect 488426 453498 488982 454054
rect 488426 417498 488982 418054
rect 488426 381498 488982 382054
rect 488426 345498 488982 346054
rect 488426 309498 488982 310054
rect 488426 273498 488982 274054
rect 488426 237498 488982 238054
rect 488426 201498 488982 202054
rect 488426 165498 488982 166054
rect 488426 129498 488982 130054
rect 488426 93498 488982 94054
rect 488426 57498 488982 58054
rect 488426 21498 488982 22054
rect 488426 -5702 488982 -5146
rect 492146 710042 492702 710598
rect 492146 673218 492702 673774
rect 492146 637218 492702 637774
rect 492146 601218 492702 601774
rect 492146 565218 492702 565774
rect 492146 529218 492702 529774
rect 492146 493218 492702 493774
rect 492146 457218 492702 457774
rect 492146 421218 492702 421774
rect 492146 385218 492702 385774
rect 492146 349218 492702 349774
rect 492146 313218 492702 313774
rect 492146 277218 492702 277774
rect 492146 241218 492702 241774
rect 492146 205218 492702 205774
rect 492146 169218 492702 169774
rect 492146 133218 492702 133774
rect 492146 97218 492702 97774
rect 492146 61218 492702 61774
rect 492146 25218 492702 25774
rect 492146 -6662 492702 -6106
rect 495866 711002 496422 711558
rect 495866 676938 496422 677494
rect 495866 640938 496422 641494
rect 495866 604938 496422 605494
rect 495866 568938 496422 569494
rect 495866 532938 496422 533494
rect 495866 496938 496422 497494
rect 495866 460938 496422 461494
rect 495866 424938 496422 425494
rect 495866 388938 496422 389494
rect 495866 352938 496422 353494
rect 495866 316938 496422 317494
rect 495866 280938 496422 281494
rect 495866 244938 496422 245494
rect 495866 208938 496422 209494
rect 495866 172938 496422 173494
rect 495866 136938 496422 137494
rect 495866 100938 496422 101494
rect 495866 64938 496422 65494
rect 495866 28938 496422 29494
rect 495866 -7622 496422 -7066
rect 505826 704282 506382 704838
rect 505826 686898 506382 687454
rect 505826 650898 506382 651454
rect 505826 614898 506382 615454
rect 505826 578898 506382 579454
rect 505826 542898 506382 543454
rect 505826 506898 506382 507454
rect 505826 470898 506382 471454
rect 505826 434898 506382 435454
rect 505826 398898 506382 399454
rect 505826 362898 506382 363454
rect 505826 326898 506382 327454
rect 505826 290898 506382 291454
rect 505826 254898 506382 255454
rect 505826 218898 506382 219454
rect 505826 182898 506382 183454
rect 505826 146898 506382 147454
rect 505826 110898 506382 111454
rect 505826 74898 506382 75454
rect 505826 38898 506382 39454
rect 505826 2898 506382 3454
rect 505826 -902 506382 -346
rect 509546 705242 510102 705798
rect 509546 690618 510102 691174
rect 509546 654618 510102 655174
rect 509546 618618 510102 619174
rect 509546 582618 510102 583174
rect 509546 546618 510102 547174
rect 509546 510618 510102 511174
rect 509546 474618 510102 475174
rect 509546 438618 510102 439174
rect 509546 402618 510102 403174
rect 509546 366618 510102 367174
rect 509546 330618 510102 331174
rect 509546 294618 510102 295174
rect 509546 258618 510102 259174
rect 509546 222618 510102 223174
rect 509546 186618 510102 187174
rect 509546 150618 510102 151174
rect 509546 114618 510102 115174
rect 509546 78618 510102 79174
rect 509546 42618 510102 43174
rect 509546 6618 510102 7174
rect 509546 -1862 510102 -1306
rect 513266 706202 513822 706758
rect 513266 694338 513822 694894
rect 513266 658338 513822 658894
rect 513266 622338 513822 622894
rect 513266 586338 513822 586894
rect 513266 550338 513822 550894
rect 513266 514338 513822 514894
rect 513266 478338 513822 478894
rect 513266 442338 513822 442894
rect 513266 406338 513822 406894
rect 513266 370338 513822 370894
rect 513266 334338 513822 334894
rect 513266 298338 513822 298894
rect 513266 262338 513822 262894
rect 513266 226338 513822 226894
rect 513266 190338 513822 190894
rect 513266 154338 513822 154894
rect 513266 118338 513822 118894
rect 513266 82338 513822 82894
rect 513266 46338 513822 46894
rect 513266 10338 513822 10894
rect 513266 -2822 513822 -2266
rect 516986 707162 517542 707718
rect 516986 698058 517542 698614
rect 516986 662058 517542 662614
rect 516986 626058 517542 626614
rect 516986 590058 517542 590614
rect 516986 554058 517542 554614
rect 516986 518058 517542 518614
rect 516986 482058 517542 482614
rect 516986 446058 517542 446614
rect 516986 410058 517542 410614
rect 516986 374058 517542 374614
rect 516986 338058 517542 338614
rect 516986 302058 517542 302614
rect 516986 266058 517542 266614
rect 516986 230058 517542 230614
rect 516986 194058 517542 194614
rect 516986 158058 517542 158614
rect 516986 122058 517542 122614
rect 516986 86058 517542 86614
rect 516986 50058 517542 50614
rect 516986 14058 517542 14614
rect 516986 -3782 517542 -3226
rect 520706 708122 521262 708678
rect 520706 665778 521262 666334
rect 520706 629778 521262 630334
rect 520706 593778 521262 594334
rect 520706 557778 521262 558334
rect 520706 521778 521262 522334
rect 520706 485778 521262 486334
rect 520706 449778 521262 450334
rect 520706 413778 521262 414334
rect 520706 377778 521262 378334
rect 520706 341778 521262 342334
rect 520706 305778 521262 306334
rect 520706 269778 521262 270334
rect 520706 233778 521262 234334
rect 520706 197778 521262 198334
rect 520706 161778 521262 162334
rect 520706 125778 521262 126334
rect 520706 89778 521262 90334
rect 520706 53778 521262 54334
rect 520706 17778 521262 18334
rect 520706 -4742 521262 -4186
rect 524426 709082 524982 709638
rect 524426 669498 524982 670054
rect 524426 633498 524982 634054
rect 524426 597498 524982 598054
rect 524426 561498 524982 562054
rect 524426 525498 524982 526054
rect 524426 489498 524982 490054
rect 524426 453498 524982 454054
rect 524426 417498 524982 418054
rect 524426 381498 524982 382054
rect 524426 345498 524982 346054
rect 524426 309498 524982 310054
rect 524426 273498 524982 274054
rect 524426 237498 524982 238054
rect 524426 201498 524982 202054
rect 524426 165498 524982 166054
rect 524426 129498 524982 130054
rect 524426 93498 524982 94054
rect 524426 57498 524982 58054
rect 524426 21498 524982 22054
rect 524426 -5702 524982 -5146
rect 528146 710042 528702 710598
rect 528146 673218 528702 673774
rect 528146 637218 528702 637774
rect 528146 601218 528702 601774
rect 528146 565218 528702 565774
rect 528146 529218 528702 529774
rect 528146 493218 528702 493774
rect 528146 457218 528702 457774
rect 528146 421218 528702 421774
rect 528146 385218 528702 385774
rect 528146 349218 528702 349774
rect 528146 313218 528702 313774
rect 528146 277218 528702 277774
rect 528146 241218 528702 241774
rect 528146 205218 528702 205774
rect 528146 169218 528702 169774
rect 528146 133218 528702 133774
rect 528146 97218 528702 97774
rect 528146 61218 528702 61774
rect 528146 25218 528702 25774
rect 528146 -6662 528702 -6106
rect 531866 711002 532422 711558
rect 531866 676938 532422 677494
rect 531866 640938 532422 641494
rect 531866 604938 532422 605494
rect 531866 568938 532422 569494
rect 531866 532938 532422 533494
rect 531866 496938 532422 497494
rect 531866 460938 532422 461494
rect 531866 424938 532422 425494
rect 531866 388938 532422 389494
rect 531866 352938 532422 353494
rect 531866 316938 532422 317494
rect 531866 280938 532422 281494
rect 531866 244938 532422 245494
rect 531866 208938 532422 209494
rect 531866 172938 532422 173494
rect 531866 136938 532422 137494
rect 531866 100938 532422 101494
rect 531866 64938 532422 65494
rect 531866 28938 532422 29494
rect 531866 -7622 532422 -7066
rect 541826 704282 542382 704838
rect 541826 686898 542382 687454
rect 541826 650898 542382 651454
rect 541826 614898 542382 615454
rect 541826 578898 542382 579454
rect 541826 542898 542382 543454
rect 541826 506898 542382 507454
rect 541826 470898 542382 471454
rect 541826 434898 542382 435454
rect 541826 398898 542382 399454
rect 541826 362898 542382 363454
rect 541826 326898 542382 327454
rect 541826 290898 542382 291454
rect 541826 254898 542382 255454
rect 541826 218898 542382 219454
rect 541826 182898 542382 183454
rect 541826 146898 542382 147454
rect 541826 110898 542382 111454
rect 541826 74898 542382 75454
rect 541826 38898 542382 39454
rect 541826 2898 542382 3454
rect 541826 -902 542382 -346
rect 545546 705242 546102 705798
rect 545546 690618 546102 691174
rect 545546 654618 546102 655174
rect 545546 618618 546102 619174
rect 545546 582618 546102 583174
rect 545546 546618 546102 547174
rect 545546 510618 546102 511174
rect 545546 474618 546102 475174
rect 545546 438618 546102 439174
rect 545546 402618 546102 403174
rect 545546 366618 546102 367174
rect 545546 330618 546102 331174
rect 545546 294618 546102 295174
rect 545546 258618 546102 259174
rect 545546 222618 546102 223174
rect 545546 186618 546102 187174
rect 545546 150618 546102 151174
rect 545546 114618 546102 115174
rect 545546 78618 546102 79174
rect 545546 42618 546102 43174
rect 545546 6618 546102 7174
rect 545546 -1862 546102 -1306
rect 549266 706202 549822 706758
rect 549266 694338 549822 694894
rect 549266 658338 549822 658894
rect 549266 622338 549822 622894
rect 549266 586338 549822 586894
rect 549266 550338 549822 550894
rect 549266 514338 549822 514894
rect 549266 478338 549822 478894
rect 549266 442338 549822 442894
rect 549266 406338 549822 406894
rect 549266 370338 549822 370894
rect 549266 334338 549822 334894
rect 549266 298338 549822 298894
rect 549266 262338 549822 262894
rect 549266 226338 549822 226894
rect 549266 190338 549822 190894
rect 549266 154338 549822 154894
rect 549266 118338 549822 118894
rect 549266 82338 549822 82894
rect 549266 46338 549822 46894
rect 549266 10338 549822 10894
rect 549266 -2822 549822 -2266
rect 552986 707162 553542 707718
rect 552986 698058 553542 698614
rect 552986 662058 553542 662614
rect 552986 626058 553542 626614
rect 552986 590058 553542 590614
rect 552986 554058 553542 554614
rect 552986 518058 553542 518614
rect 552986 482058 553542 482614
rect 552986 446058 553542 446614
rect 552986 410058 553542 410614
rect 552986 374058 553542 374614
rect 552986 338058 553542 338614
rect 552986 302058 553542 302614
rect 552986 266058 553542 266614
rect 552986 230058 553542 230614
rect 552986 194058 553542 194614
rect 552986 158058 553542 158614
rect 552986 122058 553542 122614
rect 552986 86058 553542 86614
rect 552986 50058 553542 50614
rect 552986 14058 553542 14614
rect 552986 -3782 553542 -3226
rect 556706 708122 557262 708678
rect 556706 665778 557262 666334
rect 556706 629778 557262 630334
rect 556706 593778 557262 594334
rect 556706 557778 557262 558334
rect 556706 521778 557262 522334
rect 556706 485778 557262 486334
rect 556706 449778 557262 450334
rect 556706 413778 557262 414334
rect 556706 377778 557262 378334
rect 556706 341778 557262 342334
rect 556706 305778 557262 306334
rect 556706 269778 557262 270334
rect 556706 233778 557262 234334
rect 556706 197778 557262 198334
rect 556706 161778 557262 162334
rect 556706 125778 557262 126334
rect 556706 89778 557262 90334
rect 556706 53778 557262 54334
rect 556706 17778 557262 18334
rect 556706 -4742 557262 -4186
rect 560426 709082 560982 709638
rect 560426 669498 560982 670054
rect 560426 633498 560982 634054
rect 560426 597498 560982 598054
rect 560426 561498 560982 562054
rect 560426 525498 560982 526054
rect 560426 489498 560982 490054
rect 560426 453498 560982 454054
rect 560426 417498 560982 418054
rect 560426 381498 560982 382054
rect 560426 345498 560982 346054
rect 560426 309498 560982 310054
rect 560426 273498 560982 274054
rect 560426 237498 560982 238054
rect 560426 201498 560982 202054
rect 560426 165498 560982 166054
rect 560426 129498 560982 130054
rect 560426 93498 560982 94054
rect 560426 57498 560982 58054
rect 560426 21498 560982 22054
rect 560426 -5702 560982 -5146
rect 564146 710042 564702 710598
rect 564146 673218 564702 673774
rect 564146 637218 564702 637774
rect 564146 601218 564702 601774
rect 564146 565218 564702 565774
rect 564146 529218 564702 529774
rect 564146 493218 564702 493774
rect 564146 457218 564702 457774
rect 564146 421218 564702 421774
rect 564146 385218 564702 385774
rect 564146 349218 564702 349774
rect 564146 313218 564702 313774
rect 564146 277218 564702 277774
rect 564146 241218 564702 241774
rect 564146 205218 564702 205774
rect 564146 169218 564702 169774
rect 564146 133218 564702 133774
rect 564146 97218 564702 97774
rect 564146 61218 564702 61774
rect 564146 25218 564702 25774
rect 564146 -6662 564702 -6106
rect 567866 711002 568422 711558
rect 567866 676938 568422 677494
rect 567866 640938 568422 641494
rect 567866 604938 568422 605494
rect 567866 568938 568422 569494
rect 567866 532938 568422 533494
rect 567866 496938 568422 497494
rect 567866 460938 568422 461494
rect 567866 424938 568422 425494
rect 567866 388938 568422 389494
rect 567866 352938 568422 353494
rect 567866 316938 568422 317494
rect 567866 280938 568422 281494
rect 567866 244938 568422 245494
rect 567866 208938 568422 209494
rect 567866 172938 568422 173494
rect 567866 136938 568422 137494
rect 567866 100938 568422 101494
rect 567866 64938 568422 65494
rect 567866 28938 568422 29494
rect 567866 -7622 568422 -7066
rect 577826 704282 578382 704838
rect 577826 686898 578382 687454
rect 577826 650898 578382 651454
rect 592062 711002 592618 711558
rect 591102 710042 591658 710598
rect 590142 709082 590698 709638
rect 589182 708122 589738 708678
rect 588222 707162 588778 707718
rect 587262 706202 587818 706758
rect 581546 705242 582102 705798
rect 586302 705242 586858 705798
rect 581546 690618 582102 691174
rect 581546 654618 582102 655174
rect 581546 618618 582102 619174
rect 577826 614898 578382 615454
rect 577826 578898 578382 579454
rect 577826 542898 578382 543454
rect 577826 506898 578382 507454
rect 577826 470898 578382 471454
rect 577826 434898 578382 435454
rect 577826 398898 578382 399454
rect 577826 362898 578382 363454
rect 577826 326898 578382 327454
rect 577826 290898 578382 291454
rect 577826 254898 578382 255454
rect 577826 218898 578382 219454
rect 577826 182898 578382 183454
rect 577826 146898 578382 147454
rect 577826 110898 578382 111454
rect 577826 74898 578382 75454
rect 577826 38898 578382 39454
rect 577826 2898 578382 3454
rect 581546 582618 582102 583174
rect 581546 546618 582102 547174
rect 581546 510618 582102 511174
rect 581546 474618 582102 475174
rect 581546 438618 582102 439174
rect 581546 402618 582102 403174
rect 581546 366618 582102 367174
rect 581546 330618 582102 331174
rect 581546 294618 582102 295174
rect 581546 258618 582102 259174
rect 581546 222618 582102 223174
rect 581546 186618 582102 187174
rect 581546 150618 582102 151174
rect 581546 114618 582102 115174
rect 581546 78618 582102 79174
rect 581546 42618 582102 43174
rect 581546 6618 582102 7174
rect 577826 -902 578382 -346
rect 585342 704282 585898 704838
rect 585342 686898 585898 687454
rect 585342 650898 585898 651454
rect 585342 614898 585898 615454
rect 585342 578898 585898 579454
rect 585342 542898 585898 543454
rect 585342 506898 585898 507454
rect 585342 470898 585898 471454
rect 585342 434898 585898 435454
rect 585342 398898 585898 399454
rect 585342 362898 585898 363454
rect 585342 326898 585898 327454
rect 585342 290898 585898 291454
rect 585342 254898 585898 255454
rect 585342 218898 585898 219454
rect 585342 182898 585898 183454
rect 585342 146898 585898 147454
rect 585342 110898 585898 111454
rect 585342 74898 585898 75454
rect 585342 38898 585898 39454
rect 585342 2898 585898 3454
rect 585342 -902 585898 -346
rect 586302 690618 586858 691174
rect 586302 654618 586858 655174
rect 586302 618618 586858 619174
rect 586302 582618 586858 583174
rect 586302 546618 586858 547174
rect 586302 510618 586858 511174
rect 586302 474618 586858 475174
rect 586302 438618 586858 439174
rect 586302 402618 586858 403174
rect 586302 366618 586858 367174
rect 586302 330618 586858 331174
rect 586302 294618 586858 295174
rect 586302 258618 586858 259174
rect 586302 222618 586858 223174
rect 586302 186618 586858 187174
rect 586302 150618 586858 151174
rect 586302 114618 586858 115174
rect 586302 78618 586858 79174
rect 586302 42618 586858 43174
rect 586302 6618 586858 7174
rect 581546 -1862 582102 -1306
rect 586302 -1862 586858 -1306
rect 587262 694338 587818 694894
rect 587262 658338 587818 658894
rect 587262 622338 587818 622894
rect 587262 586338 587818 586894
rect 587262 550338 587818 550894
rect 587262 514338 587818 514894
rect 587262 478338 587818 478894
rect 587262 442338 587818 442894
rect 587262 406338 587818 406894
rect 587262 370338 587818 370894
rect 587262 334338 587818 334894
rect 587262 298338 587818 298894
rect 587262 262338 587818 262894
rect 587262 226338 587818 226894
rect 587262 190338 587818 190894
rect 587262 154338 587818 154894
rect 587262 118338 587818 118894
rect 587262 82338 587818 82894
rect 587262 46338 587818 46894
rect 587262 10338 587818 10894
rect 587262 -2822 587818 -2266
rect 588222 698058 588778 698614
rect 588222 662058 588778 662614
rect 588222 626058 588778 626614
rect 588222 590058 588778 590614
rect 588222 554058 588778 554614
rect 588222 518058 588778 518614
rect 588222 482058 588778 482614
rect 588222 446058 588778 446614
rect 588222 410058 588778 410614
rect 588222 374058 588778 374614
rect 588222 338058 588778 338614
rect 588222 302058 588778 302614
rect 588222 266058 588778 266614
rect 588222 230058 588778 230614
rect 588222 194058 588778 194614
rect 588222 158058 588778 158614
rect 588222 122058 588778 122614
rect 588222 86058 588778 86614
rect 588222 50058 588778 50614
rect 588222 14058 588778 14614
rect 588222 -3782 588778 -3226
rect 589182 665778 589738 666334
rect 589182 629778 589738 630334
rect 589182 593778 589738 594334
rect 589182 557778 589738 558334
rect 589182 521778 589738 522334
rect 589182 485778 589738 486334
rect 589182 449778 589738 450334
rect 589182 413778 589738 414334
rect 589182 377778 589738 378334
rect 589182 341778 589738 342334
rect 589182 305778 589738 306334
rect 589182 269778 589738 270334
rect 589182 233778 589738 234334
rect 589182 197778 589738 198334
rect 589182 161778 589738 162334
rect 589182 125778 589738 126334
rect 589182 89778 589738 90334
rect 589182 53778 589738 54334
rect 589182 17778 589738 18334
rect 589182 -4742 589738 -4186
rect 590142 669498 590698 670054
rect 590142 633498 590698 634054
rect 590142 597498 590698 598054
rect 590142 561498 590698 562054
rect 590142 525498 590698 526054
rect 590142 489498 590698 490054
rect 590142 453498 590698 454054
rect 590142 417498 590698 418054
rect 590142 381498 590698 382054
rect 590142 345498 590698 346054
rect 590142 309498 590698 310054
rect 590142 273498 590698 274054
rect 590142 237498 590698 238054
rect 590142 201498 590698 202054
rect 590142 165498 590698 166054
rect 590142 129498 590698 130054
rect 590142 93498 590698 94054
rect 590142 57498 590698 58054
rect 590142 21498 590698 22054
rect 590142 -5702 590698 -5146
rect 591102 673218 591658 673774
rect 591102 637218 591658 637774
rect 591102 601218 591658 601774
rect 591102 565218 591658 565774
rect 591102 529218 591658 529774
rect 591102 493218 591658 493774
rect 591102 457218 591658 457774
rect 591102 421218 591658 421774
rect 591102 385218 591658 385774
rect 591102 349218 591658 349774
rect 591102 313218 591658 313774
rect 591102 277218 591658 277774
rect 591102 241218 591658 241774
rect 591102 205218 591658 205774
rect 591102 169218 591658 169774
rect 591102 133218 591658 133774
rect 591102 97218 591658 97774
rect 591102 61218 591658 61774
rect 591102 25218 591658 25774
rect 591102 -6662 591658 -6106
rect 592062 676938 592618 677494
rect 592062 640938 592618 641494
rect 592062 604938 592618 605494
rect 592062 568938 592618 569494
rect 592062 532938 592618 533494
rect 592062 496938 592618 497494
rect 592062 460938 592618 461494
rect 592062 424938 592618 425494
rect 592062 388938 592618 389494
rect 592062 352938 592618 353494
rect 592062 316938 592618 317494
rect 592062 280938 592618 281494
rect 592062 244938 592618 245494
rect 592062 208938 592618 209494
rect 592062 172938 592618 173494
rect 592062 136938 592618 137494
rect 592062 100938 592618 101494
rect 592062 64938 592618 65494
rect 592062 28938 592618 29494
rect 592062 -7622 592618 -7066
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711002 -8694 711558
rect -8138 711002 27866 711558
rect 28422 711002 63866 711558
rect 64422 711002 99866 711558
rect 100422 711002 135866 711558
rect 136422 711002 171866 711558
rect 172422 711002 207866 711558
rect 208422 711002 243866 711558
rect 244422 711002 279866 711558
rect 280422 711002 315866 711558
rect 316422 711002 351866 711558
rect 352422 711002 387866 711558
rect 388422 711002 423866 711558
rect 424422 711002 459866 711558
rect 460422 711002 495866 711558
rect 496422 711002 531866 711558
rect 532422 711002 567866 711558
rect 568422 711002 592062 711558
rect 592618 711002 592650 711558
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710042 -7734 710598
rect -7178 710042 24146 710598
rect 24702 710042 60146 710598
rect 60702 710042 96146 710598
rect 96702 710042 132146 710598
rect 132702 710042 168146 710598
rect 168702 710042 204146 710598
rect 204702 710042 240146 710598
rect 240702 710042 276146 710598
rect 276702 710042 312146 710598
rect 312702 710042 348146 710598
rect 348702 710042 384146 710598
rect 384702 710042 420146 710598
rect 420702 710042 456146 710598
rect 456702 710042 492146 710598
rect 492702 710042 528146 710598
rect 528702 710042 564146 710598
rect 564702 710042 591102 710598
rect 591658 710042 591690 710598
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709082 -6774 709638
rect -6218 709082 20426 709638
rect 20982 709082 56426 709638
rect 56982 709082 92426 709638
rect 92982 709082 128426 709638
rect 128982 709082 164426 709638
rect 164982 709082 200426 709638
rect 200982 709082 236426 709638
rect 236982 709082 272426 709638
rect 272982 709082 308426 709638
rect 308982 709082 344426 709638
rect 344982 709082 380426 709638
rect 380982 709082 416426 709638
rect 416982 709082 452426 709638
rect 452982 709082 488426 709638
rect 488982 709082 524426 709638
rect 524982 709082 560426 709638
rect 560982 709082 590142 709638
rect 590698 709082 590730 709638
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708122 -5814 708678
rect -5258 708122 16706 708678
rect 17262 708122 52706 708678
rect 53262 708122 88706 708678
rect 89262 708122 124706 708678
rect 125262 708122 160706 708678
rect 161262 708122 196706 708678
rect 197262 708122 232706 708678
rect 233262 708122 268706 708678
rect 269262 708122 304706 708678
rect 305262 708122 340706 708678
rect 341262 708122 376706 708678
rect 377262 708122 412706 708678
rect 413262 708122 448706 708678
rect 449262 708122 484706 708678
rect 485262 708122 520706 708678
rect 521262 708122 556706 708678
rect 557262 708122 589182 708678
rect 589738 708122 589770 708678
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707162 -4854 707718
rect -4298 707162 12986 707718
rect 13542 707162 48986 707718
rect 49542 707162 84986 707718
rect 85542 707162 120986 707718
rect 121542 707162 156986 707718
rect 157542 707162 192986 707718
rect 193542 707162 228986 707718
rect 229542 707162 264986 707718
rect 265542 707162 300986 707718
rect 301542 707162 336986 707718
rect 337542 707162 372986 707718
rect 373542 707162 408986 707718
rect 409542 707162 444986 707718
rect 445542 707162 480986 707718
rect 481542 707162 516986 707718
rect 517542 707162 552986 707718
rect 553542 707162 588222 707718
rect 588778 707162 588810 707718
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706202 -3894 706758
rect -3338 706202 9266 706758
rect 9822 706202 45266 706758
rect 45822 706202 81266 706758
rect 81822 706202 117266 706758
rect 117822 706202 153266 706758
rect 153822 706202 189266 706758
rect 189822 706202 225266 706758
rect 225822 706202 261266 706758
rect 261822 706202 297266 706758
rect 297822 706202 333266 706758
rect 333822 706202 369266 706758
rect 369822 706202 405266 706758
rect 405822 706202 441266 706758
rect 441822 706202 477266 706758
rect 477822 706202 513266 706758
rect 513822 706202 549266 706758
rect 549822 706202 587262 706758
rect 587818 706202 587850 706758
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705242 -2934 705798
rect -2378 705242 5546 705798
rect 6102 705242 41546 705798
rect 42102 705242 77546 705798
rect 78102 705242 113546 705798
rect 114102 705242 149546 705798
rect 150102 705242 185546 705798
rect 186102 705242 221546 705798
rect 222102 705242 257546 705798
rect 258102 705242 293546 705798
rect 294102 705242 329546 705798
rect 330102 705242 365546 705798
rect 366102 705242 401546 705798
rect 402102 705242 437546 705798
rect 438102 705242 473546 705798
rect 474102 705242 509546 705798
rect 510102 705242 545546 705798
rect 546102 705242 581546 705798
rect 582102 705242 586302 705798
rect 586858 705242 586890 705798
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704282 -1974 704838
rect -1418 704282 1826 704838
rect 2382 704282 37826 704838
rect 38382 704282 73826 704838
rect 74382 704282 109826 704838
rect 110382 704282 145826 704838
rect 146382 704282 181826 704838
rect 182382 704282 217826 704838
rect 218382 704282 253826 704838
rect 254382 704282 289826 704838
rect 290382 704282 325826 704838
rect 326382 704282 361826 704838
rect 362382 704282 397826 704838
rect 398382 704282 433826 704838
rect 434382 704282 469826 704838
rect 470382 704282 505826 704838
rect 506382 704282 541826 704838
rect 542382 704282 577826 704838
rect 578382 704282 585342 704838
rect 585898 704282 585930 704838
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698058 -4854 698614
rect -4298 698058 12986 698614
rect 13542 698058 48986 698614
rect 49542 698058 84986 698614
rect 85542 698058 120986 698614
rect 121542 698058 156986 698614
rect 157542 698058 192986 698614
rect 193542 698058 228986 698614
rect 229542 698058 264986 698614
rect 265542 698058 300986 698614
rect 301542 698058 336986 698614
rect 337542 698058 372986 698614
rect 373542 698058 408986 698614
rect 409542 698058 444986 698614
rect 445542 698058 480986 698614
rect 481542 698058 516986 698614
rect 517542 698058 552986 698614
rect 553542 698058 588222 698614
rect 588778 698058 592650 698614
rect -8726 698026 592650 698058
rect -8726 694894 592650 694926
rect -8726 694338 -3894 694894
rect -3338 694338 9266 694894
rect 9822 694338 45266 694894
rect 45822 694338 81266 694894
rect 81822 694338 117266 694894
rect 117822 694338 153266 694894
rect 153822 694338 189266 694894
rect 189822 694338 225266 694894
rect 225822 694338 261266 694894
rect 261822 694338 297266 694894
rect 297822 694338 333266 694894
rect 333822 694338 369266 694894
rect 369822 694338 405266 694894
rect 405822 694338 441266 694894
rect 441822 694338 477266 694894
rect 477822 694338 513266 694894
rect 513822 694338 549266 694894
rect 549822 694338 587262 694894
rect 587818 694338 592650 694894
rect -8726 694306 592650 694338
rect -8726 691174 592650 691206
rect -8726 690618 -2934 691174
rect -2378 690618 5546 691174
rect 6102 690618 41546 691174
rect 42102 690618 77546 691174
rect 78102 690618 113546 691174
rect 114102 690618 149546 691174
rect 150102 690618 185546 691174
rect 186102 690618 221546 691174
rect 222102 690618 257546 691174
rect 258102 690618 293546 691174
rect 294102 690618 329546 691174
rect 330102 690618 365546 691174
rect 366102 690618 401546 691174
rect 402102 690618 437546 691174
rect 438102 690618 473546 691174
rect 474102 690618 509546 691174
rect 510102 690618 545546 691174
rect 546102 690618 581546 691174
rect 582102 690618 586302 691174
rect 586858 690618 592650 691174
rect -8726 690586 592650 690618
rect -8726 687454 592650 687486
rect -8726 686898 -1974 687454
rect -1418 686898 1826 687454
rect 2382 686898 37826 687454
rect 38382 686898 73826 687454
rect 74382 686898 109826 687454
rect 110382 686898 145826 687454
rect 146382 686898 181826 687454
rect 182382 686898 217826 687454
rect 218382 686898 253826 687454
rect 254382 686898 289826 687454
rect 290382 686898 325826 687454
rect 326382 686898 361826 687454
rect 362382 686898 397826 687454
rect 398382 686898 433826 687454
rect 434382 686898 469826 687454
rect 470382 686898 505826 687454
rect 506382 686898 541826 687454
rect 542382 686898 577826 687454
rect 578382 686898 585342 687454
rect 585898 686898 592650 687454
rect -8726 686866 592650 686898
rect -8726 677494 592650 677526
rect -8726 676938 -8694 677494
rect -8138 676938 27866 677494
rect 28422 676938 63866 677494
rect 64422 676938 99866 677494
rect 100422 676938 135866 677494
rect 136422 676938 171866 677494
rect 172422 676938 207866 677494
rect 208422 676938 243866 677494
rect 244422 676938 279866 677494
rect 280422 676938 315866 677494
rect 316422 676938 351866 677494
rect 352422 676938 387866 677494
rect 388422 676938 423866 677494
rect 424422 676938 459866 677494
rect 460422 676938 495866 677494
rect 496422 676938 531866 677494
rect 532422 676938 567866 677494
rect 568422 676938 592062 677494
rect 592618 676938 592650 677494
rect -8726 676906 592650 676938
rect -8726 673774 592650 673806
rect -8726 673218 -7734 673774
rect -7178 673218 24146 673774
rect 24702 673218 60146 673774
rect 60702 673218 96146 673774
rect 96702 673218 132146 673774
rect 132702 673218 168146 673774
rect 168702 673218 204146 673774
rect 204702 673218 240146 673774
rect 240702 673218 276146 673774
rect 276702 673218 312146 673774
rect 312702 673218 348146 673774
rect 348702 673218 384146 673774
rect 384702 673218 420146 673774
rect 420702 673218 456146 673774
rect 456702 673218 492146 673774
rect 492702 673218 528146 673774
rect 528702 673218 564146 673774
rect 564702 673218 591102 673774
rect 591658 673218 592650 673774
rect -8726 673186 592650 673218
rect -8726 670054 592650 670086
rect -8726 669498 -6774 670054
rect -6218 669498 20426 670054
rect 20982 669498 56426 670054
rect 56982 669498 92426 670054
rect 92982 669498 128426 670054
rect 128982 669498 164426 670054
rect 164982 669498 200426 670054
rect 200982 669498 236426 670054
rect 236982 669498 272426 670054
rect 272982 669498 308426 670054
rect 308982 669498 344426 670054
rect 344982 669498 380426 670054
rect 380982 669498 416426 670054
rect 416982 669498 452426 670054
rect 452982 669498 488426 670054
rect 488982 669498 524426 670054
rect 524982 669498 560426 670054
rect 560982 669498 590142 670054
rect 590698 669498 592650 670054
rect -8726 669466 592650 669498
rect -8726 666334 592650 666366
rect -8726 665778 -5814 666334
rect -5258 665778 16706 666334
rect 17262 665778 52706 666334
rect 53262 665778 88706 666334
rect 89262 665778 124706 666334
rect 125262 665778 160706 666334
rect 161262 665778 196706 666334
rect 197262 665778 232706 666334
rect 233262 665778 268706 666334
rect 269262 665778 304706 666334
rect 305262 665778 340706 666334
rect 341262 665778 376706 666334
rect 377262 665778 412706 666334
rect 413262 665778 448706 666334
rect 449262 665778 484706 666334
rect 485262 665778 520706 666334
rect 521262 665778 556706 666334
rect 557262 665778 589182 666334
rect 589738 665778 592650 666334
rect -8726 665746 592650 665778
rect -8726 662614 592650 662646
rect -8726 662058 -4854 662614
rect -4298 662058 12986 662614
rect 13542 662058 48986 662614
rect 49542 662058 84986 662614
rect 85542 662058 120986 662614
rect 121542 662058 156986 662614
rect 157542 662058 192986 662614
rect 193542 662058 228986 662614
rect 229542 662058 264986 662614
rect 265542 662058 300986 662614
rect 301542 662058 336986 662614
rect 337542 662058 372986 662614
rect 373542 662058 408986 662614
rect 409542 662058 444986 662614
rect 445542 662058 480986 662614
rect 481542 662058 516986 662614
rect 517542 662058 552986 662614
rect 553542 662058 588222 662614
rect 588778 662058 592650 662614
rect -8726 662026 592650 662058
rect -8726 658894 592650 658926
rect -8726 658338 -3894 658894
rect -3338 658338 9266 658894
rect 9822 658338 45266 658894
rect 45822 658338 81266 658894
rect 81822 658338 117266 658894
rect 117822 658338 153266 658894
rect 153822 658338 189266 658894
rect 189822 658338 225266 658894
rect 225822 658338 261266 658894
rect 261822 658338 297266 658894
rect 297822 658338 333266 658894
rect 333822 658338 369266 658894
rect 369822 658338 405266 658894
rect 405822 658338 441266 658894
rect 441822 658338 477266 658894
rect 477822 658338 513266 658894
rect 513822 658338 549266 658894
rect 549822 658338 587262 658894
rect 587818 658338 592650 658894
rect -8726 658306 592650 658338
rect -8726 655174 592650 655206
rect -8726 654618 -2934 655174
rect -2378 654618 5546 655174
rect 6102 654618 41546 655174
rect 42102 654618 77546 655174
rect 78102 654618 113546 655174
rect 114102 654618 149546 655174
rect 150102 654618 185546 655174
rect 186102 654618 221546 655174
rect 222102 654618 257546 655174
rect 258102 654618 293546 655174
rect 294102 654618 329546 655174
rect 330102 654618 365546 655174
rect 366102 654618 401546 655174
rect 402102 654618 437546 655174
rect 438102 654618 473546 655174
rect 474102 654618 509546 655174
rect 510102 654618 545546 655174
rect 546102 654618 581546 655174
rect 582102 654618 586302 655174
rect 586858 654618 592650 655174
rect -8726 654586 592650 654618
rect -8726 651454 592650 651486
rect -8726 650898 -1974 651454
rect -1418 650898 1826 651454
rect 2382 650898 37826 651454
rect 38382 650898 73826 651454
rect 74382 650898 109826 651454
rect 110382 650898 145826 651454
rect 146382 650898 181826 651454
rect 182382 650898 217826 651454
rect 218382 650898 253826 651454
rect 254382 650898 289826 651454
rect 290382 650898 325826 651454
rect 326382 650898 361826 651454
rect 362382 650898 397826 651454
rect 398382 650898 433826 651454
rect 434382 650898 469826 651454
rect 470382 650898 505826 651454
rect 506382 650898 541826 651454
rect 542382 650898 577826 651454
rect 578382 650898 585342 651454
rect 585898 650898 592650 651454
rect -8726 650866 592650 650898
rect -8726 641494 592650 641526
rect -8726 640938 -8694 641494
rect -8138 640938 27866 641494
rect 28422 640938 63866 641494
rect 64422 640938 99866 641494
rect 100422 640938 135866 641494
rect 136422 640938 171866 641494
rect 172422 640938 207866 641494
rect 208422 640938 243866 641494
rect 244422 640938 279866 641494
rect 280422 640938 315866 641494
rect 316422 640938 351866 641494
rect 352422 640938 387866 641494
rect 388422 640938 423866 641494
rect 424422 640938 459866 641494
rect 460422 640938 495866 641494
rect 496422 640938 531866 641494
rect 532422 640938 567866 641494
rect 568422 640938 592062 641494
rect 592618 640938 592650 641494
rect -8726 640906 592650 640938
rect -8726 637774 592650 637806
rect -8726 637218 -7734 637774
rect -7178 637218 24146 637774
rect 24702 637218 60146 637774
rect 60702 637218 96146 637774
rect 96702 637218 132146 637774
rect 132702 637218 168146 637774
rect 168702 637218 204146 637774
rect 204702 637218 240146 637774
rect 240702 637218 276146 637774
rect 276702 637218 312146 637774
rect 312702 637218 348146 637774
rect 348702 637218 384146 637774
rect 384702 637218 420146 637774
rect 420702 637218 456146 637774
rect 456702 637218 492146 637774
rect 492702 637218 528146 637774
rect 528702 637218 564146 637774
rect 564702 637218 591102 637774
rect 591658 637218 592650 637774
rect -8726 637186 592650 637218
rect -8726 634054 592650 634086
rect -8726 633498 -6774 634054
rect -6218 633498 20426 634054
rect 20982 633498 56426 634054
rect 56982 633498 92426 634054
rect 92982 633498 128426 634054
rect 128982 633498 164426 634054
rect 164982 633498 200426 634054
rect 200982 633498 236426 634054
rect 236982 633498 272426 634054
rect 272982 633498 308426 634054
rect 308982 633498 344426 634054
rect 344982 633498 380426 634054
rect 380982 633498 416426 634054
rect 416982 633498 452426 634054
rect 452982 633498 488426 634054
rect 488982 633498 524426 634054
rect 524982 633498 560426 634054
rect 560982 633498 590142 634054
rect 590698 633498 592650 634054
rect -8726 633466 592650 633498
rect -8726 630334 592650 630366
rect -8726 629778 -5814 630334
rect -5258 629778 16706 630334
rect 17262 629778 52706 630334
rect 53262 629778 88706 630334
rect 89262 629778 124706 630334
rect 125262 629778 160706 630334
rect 161262 629778 196706 630334
rect 197262 629778 232706 630334
rect 233262 629778 268706 630334
rect 269262 629778 304706 630334
rect 305262 629778 340706 630334
rect 341262 629778 376706 630334
rect 377262 629778 412706 630334
rect 413262 629778 448706 630334
rect 449262 629778 484706 630334
rect 485262 629778 520706 630334
rect 521262 629778 556706 630334
rect 557262 629778 589182 630334
rect 589738 629778 592650 630334
rect -8726 629746 592650 629778
rect -8726 626614 592650 626646
rect -8726 626058 -4854 626614
rect -4298 626058 12986 626614
rect 13542 626058 48986 626614
rect 49542 626058 84986 626614
rect 85542 626058 120986 626614
rect 121542 626058 156986 626614
rect 157542 626058 192986 626614
rect 193542 626058 228986 626614
rect 229542 626058 264986 626614
rect 265542 626058 300986 626614
rect 301542 626058 336986 626614
rect 337542 626058 372986 626614
rect 373542 626058 408986 626614
rect 409542 626058 444986 626614
rect 445542 626058 480986 626614
rect 481542 626058 516986 626614
rect 517542 626058 552986 626614
rect 553542 626058 588222 626614
rect 588778 626058 592650 626614
rect -8726 626026 592650 626058
rect -8726 622894 592650 622926
rect -8726 622338 -3894 622894
rect -3338 622338 9266 622894
rect 9822 622338 45266 622894
rect 45822 622338 81266 622894
rect 81822 622338 117266 622894
rect 117822 622338 153266 622894
rect 153822 622338 189266 622894
rect 189822 622338 225266 622894
rect 225822 622338 261266 622894
rect 261822 622338 297266 622894
rect 297822 622338 333266 622894
rect 333822 622338 369266 622894
rect 369822 622338 405266 622894
rect 405822 622338 441266 622894
rect 441822 622338 477266 622894
rect 477822 622338 513266 622894
rect 513822 622338 549266 622894
rect 549822 622338 587262 622894
rect 587818 622338 592650 622894
rect -8726 622306 592650 622338
rect -8726 619174 592650 619206
rect -8726 618618 -2934 619174
rect -2378 618618 5546 619174
rect 6102 618618 41546 619174
rect 42102 618618 77546 619174
rect 78102 618618 113546 619174
rect 114102 618618 149546 619174
rect 150102 618618 185546 619174
rect 186102 618618 221546 619174
rect 222102 618618 257546 619174
rect 258102 618618 293546 619174
rect 294102 618618 329546 619174
rect 330102 618618 365546 619174
rect 366102 618618 401546 619174
rect 402102 618618 437546 619174
rect 438102 618618 473546 619174
rect 474102 618618 509546 619174
rect 510102 618618 545546 619174
rect 546102 618618 581546 619174
rect 582102 618618 586302 619174
rect 586858 618618 592650 619174
rect -8726 618586 592650 618618
rect -8726 615454 592650 615486
rect -8726 614898 -1974 615454
rect -1418 614898 1826 615454
rect 2382 614898 37826 615454
rect 38382 614898 73826 615454
rect 74382 614898 109826 615454
rect 110382 614898 145826 615454
rect 146382 614898 181826 615454
rect 182382 614898 217826 615454
rect 218382 614898 253826 615454
rect 254382 614898 289826 615454
rect 290382 614898 325826 615454
rect 326382 614898 361826 615454
rect 362382 614898 397826 615454
rect 398382 614898 433826 615454
rect 434382 614898 469826 615454
rect 470382 614898 505826 615454
rect 506382 614898 541826 615454
rect 542382 614898 577826 615454
rect 578382 614898 585342 615454
rect 585898 614898 592650 615454
rect -8726 614866 592650 614898
rect -8726 605494 592650 605526
rect -8726 604938 -8694 605494
rect -8138 604938 27866 605494
rect 28422 604938 63866 605494
rect 64422 604938 99866 605494
rect 100422 604938 135866 605494
rect 136422 604938 171866 605494
rect 172422 604938 207866 605494
rect 208422 604938 243866 605494
rect 244422 604938 279866 605494
rect 280422 604938 315866 605494
rect 316422 604938 351866 605494
rect 352422 604938 387866 605494
rect 388422 604938 423866 605494
rect 424422 604938 459866 605494
rect 460422 604938 495866 605494
rect 496422 604938 531866 605494
rect 532422 604938 567866 605494
rect 568422 604938 592062 605494
rect 592618 604938 592650 605494
rect -8726 604906 592650 604938
rect -8726 601774 592650 601806
rect -8726 601218 -7734 601774
rect -7178 601218 24146 601774
rect 24702 601218 60146 601774
rect 60702 601218 96146 601774
rect 96702 601218 132146 601774
rect 132702 601218 168146 601774
rect 168702 601218 204146 601774
rect 204702 601218 240146 601774
rect 240702 601218 276146 601774
rect 276702 601218 312146 601774
rect 312702 601218 348146 601774
rect 348702 601218 384146 601774
rect 384702 601218 420146 601774
rect 420702 601218 456146 601774
rect 456702 601218 492146 601774
rect 492702 601218 528146 601774
rect 528702 601218 564146 601774
rect 564702 601218 591102 601774
rect 591658 601218 592650 601774
rect -8726 601186 592650 601218
rect -8726 598054 592650 598086
rect -8726 597498 -6774 598054
rect -6218 597498 20426 598054
rect 20982 597498 56426 598054
rect 56982 597498 92426 598054
rect 92982 597498 128426 598054
rect 128982 597498 164426 598054
rect 164982 597498 200426 598054
rect 200982 597498 236426 598054
rect 236982 597498 272426 598054
rect 272982 597498 308426 598054
rect 308982 597498 344426 598054
rect 344982 597498 380426 598054
rect 380982 597498 416426 598054
rect 416982 597498 452426 598054
rect 452982 597498 488426 598054
rect 488982 597498 524426 598054
rect 524982 597498 560426 598054
rect 560982 597498 590142 598054
rect 590698 597498 592650 598054
rect -8726 597466 592650 597498
rect -8726 594334 592650 594366
rect -8726 593778 -5814 594334
rect -5258 593778 16706 594334
rect 17262 593778 52706 594334
rect 53262 593778 88706 594334
rect 89262 593778 124706 594334
rect 125262 593778 160706 594334
rect 161262 593778 196706 594334
rect 197262 593778 232706 594334
rect 233262 593778 268706 594334
rect 269262 593778 304706 594334
rect 305262 593778 340706 594334
rect 341262 593778 376706 594334
rect 377262 593778 412706 594334
rect 413262 593778 448706 594334
rect 449262 593778 484706 594334
rect 485262 593778 520706 594334
rect 521262 593778 556706 594334
rect 557262 593778 589182 594334
rect 589738 593778 592650 594334
rect -8726 593746 592650 593778
rect -8726 590614 592650 590646
rect -8726 590058 -4854 590614
rect -4298 590058 12986 590614
rect 13542 590058 48986 590614
rect 49542 590058 84986 590614
rect 85542 590058 120986 590614
rect 121542 590058 156986 590614
rect 157542 590058 192986 590614
rect 193542 590058 228986 590614
rect 229542 590058 264986 590614
rect 265542 590058 300986 590614
rect 301542 590058 336986 590614
rect 337542 590058 372986 590614
rect 373542 590058 408986 590614
rect 409542 590058 444986 590614
rect 445542 590058 480986 590614
rect 481542 590058 516986 590614
rect 517542 590058 552986 590614
rect 553542 590058 588222 590614
rect 588778 590058 592650 590614
rect -8726 590026 592650 590058
rect -8726 586894 592650 586926
rect -8726 586338 -3894 586894
rect -3338 586338 9266 586894
rect 9822 586338 45266 586894
rect 45822 586338 81266 586894
rect 81822 586338 117266 586894
rect 117822 586338 153266 586894
rect 153822 586338 189266 586894
rect 189822 586338 225266 586894
rect 225822 586338 261266 586894
rect 261822 586338 297266 586894
rect 297822 586338 333266 586894
rect 333822 586338 369266 586894
rect 369822 586338 405266 586894
rect 405822 586338 441266 586894
rect 441822 586338 477266 586894
rect 477822 586338 513266 586894
rect 513822 586338 549266 586894
rect 549822 586338 587262 586894
rect 587818 586338 592650 586894
rect -8726 586306 592650 586338
rect -8726 583174 592650 583206
rect -8726 582618 -2934 583174
rect -2378 582618 5546 583174
rect 6102 582618 41546 583174
rect 42102 582618 77546 583174
rect 78102 582618 113546 583174
rect 114102 582618 149546 583174
rect 150102 582618 185546 583174
rect 186102 582618 221546 583174
rect 222102 582618 257546 583174
rect 258102 582618 293546 583174
rect 294102 582618 329546 583174
rect 330102 582618 365546 583174
rect 366102 582618 401546 583174
rect 402102 582618 437546 583174
rect 438102 582618 473546 583174
rect 474102 582618 509546 583174
rect 510102 582618 545546 583174
rect 546102 582618 581546 583174
rect 582102 582618 586302 583174
rect 586858 582618 592650 583174
rect -8726 582586 592650 582618
rect -8726 579454 592650 579486
rect -8726 578898 -1974 579454
rect -1418 578898 1826 579454
rect 2382 578898 37826 579454
rect 38382 578898 73826 579454
rect 74382 578898 109826 579454
rect 110382 578898 145826 579454
rect 146382 578898 181826 579454
rect 182382 578898 217826 579454
rect 218382 578898 253826 579454
rect 254382 578898 289826 579454
rect 290382 578898 325826 579454
rect 326382 578898 361826 579454
rect 362382 578898 397826 579454
rect 398382 578898 433826 579454
rect 434382 578898 469826 579454
rect 470382 578898 505826 579454
rect 506382 578898 541826 579454
rect 542382 578898 577826 579454
rect 578382 578898 585342 579454
rect 585898 578898 592650 579454
rect -8726 578866 592650 578898
rect -8726 569494 592650 569526
rect -8726 568938 -8694 569494
rect -8138 568938 27866 569494
rect 28422 568938 63866 569494
rect 64422 568938 99866 569494
rect 100422 568938 135866 569494
rect 136422 568938 171866 569494
rect 172422 568938 207866 569494
rect 208422 568938 243866 569494
rect 244422 568938 279866 569494
rect 280422 568938 315866 569494
rect 316422 568938 351866 569494
rect 352422 568938 387866 569494
rect 388422 568938 423866 569494
rect 424422 568938 459866 569494
rect 460422 568938 495866 569494
rect 496422 568938 531866 569494
rect 532422 568938 567866 569494
rect 568422 568938 592062 569494
rect 592618 568938 592650 569494
rect -8726 568906 592650 568938
rect -8726 565774 592650 565806
rect -8726 565218 -7734 565774
rect -7178 565218 24146 565774
rect 24702 565218 60146 565774
rect 60702 565218 96146 565774
rect 96702 565218 132146 565774
rect 132702 565218 168146 565774
rect 168702 565218 204146 565774
rect 204702 565218 240146 565774
rect 240702 565218 276146 565774
rect 276702 565218 312146 565774
rect 312702 565218 348146 565774
rect 348702 565218 384146 565774
rect 384702 565218 420146 565774
rect 420702 565218 456146 565774
rect 456702 565218 492146 565774
rect 492702 565218 528146 565774
rect 528702 565218 564146 565774
rect 564702 565218 591102 565774
rect 591658 565218 592650 565774
rect -8726 565186 592650 565218
rect -8726 562054 592650 562086
rect -8726 561498 -6774 562054
rect -6218 561498 20426 562054
rect 20982 561498 56426 562054
rect 56982 561498 92426 562054
rect 92982 561498 128426 562054
rect 128982 561498 164426 562054
rect 164982 561498 200426 562054
rect 200982 561498 236426 562054
rect 236982 561498 272426 562054
rect 272982 561498 308426 562054
rect 308982 561498 344426 562054
rect 344982 561498 380426 562054
rect 380982 561498 416426 562054
rect 416982 561498 452426 562054
rect 452982 561498 488426 562054
rect 488982 561498 524426 562054
rect 524982 561498 560426 562054
rect 560982 561498 590142 562054
rect 590698 561498 592650 562054
rect -8726 561466 592650 561498
rect -8726 558334 592650 558366
rect -8726 557778 -5814 558334
rect -5258 557778 16706 558334
rect 17262 557778 52706 558334
rect 53262 557778 88706 558334
rect 89262 557778 124706 558334
rect 125262 557778 160706 558334
rect 161262 557778 196706 558334
rect 197262 557778 232706 558334
rect 233262 557778 268706 558334
rect 269262 557778 304706 558334
rect 305262 557778 340706 558334
rect 341262 557778 376706 558334
rect 377262 557778 412706 558334
rect 413262 557778 448706 558334
rect 449262 557778 484706 558334
rect 485262 557778 520706 558334
rect 521262 557778 556706 558334
rect 557262 557778 589182 558334
rect 589738 557778 592650 558334
rect -8726 557746 592650 557778
rect -8726 554614 592650 554646
rect -8726 554058 -4854 554614
rect -4298 554058 12986 554614
rect 13542 554058 48986 554614
rect 49542 554058 84986 554614
rect 85542 554058 120986 554614
rect 121542 554058 156986 554614
rect 157542 554058 192986 554614
rect 193542 554058 228986 554614
rect 229542 554058 264986 554614
rect 265542 554058 300986 554614
rect 301542 554058 336986 554614
rect 337542 554058 372986 554614
rect 373542 554058 408986 554614
rect 409542 554058 444986 554614
rect 445542 554058 480986 554614
rect 481542 554058 516986 554614
rect 517542 554058 552986 554614
rect 553542 554058 588222 554614
rect 588778 554058 592650 554614
rect -8726 554026 592650 554058
rect -8726 550894 592650 550926
rect -8726 550338 -3894 550894
rect -3338 550338 9266 550894
rect 9822 550338 45266 550894
rect 45822 550338 81266 550894
rect 81822 550338 117266 550894
rect 117822 550338 153266 550894
rect 153822 550338 189266 550894
rect 189822 550338 225266 550894
rect 225822 550338 261266 550894
rect 261822 550338 297266 550894
rect 297822 550338 333266 550894
rect 333822 550338 369266 550894
rect 369822 550338 405266 550894
rect 405822 550338 441266 550894
rect 441822 550338 477266 550894
rect 477822 550338 513266 550894
rect 513822 550338 549266 550894
rect 549822 550338 587262 550894
rect 587818 550338 592650 550894
rect -8726 550306 592650 550338
rect -8726 547174 592650 547206
rect -8726 546618 -2934 547174
rect -2378 546618 5546 547174
rect 6102 546618 41546 547174
rect 42102 546618 77546 547174
rect 78102 546618 113546 547174
rect 114102 546618 149546 547174
rect 150102 546618 185546 547174
rect 186102 546618 221546 547174
rect 222102 546618 257546 547174
rect 258102 546618 293546 547174
rect 294102 546618 329546 547174
rect 330102 546618 365546 547174
rect 366102 546618 401546 547174
rect 402102 546618 437546 547174
rect 438102 546618 473546 547174
rect 474102 546618 509546 547174
rect 510102 546618 545546 547174
rect 546102 546618 581546 547174
rect 582102 546618 586302 547174
rect 586858 546618 592650 547174
rect -8726 546586 592650 546618
rect -8726 543454 592650 543486
rect -8726 542898 -1974 543454
rect -1418 542898 1826 543454
rect 2382 542898 37826 543454
rect 38382 542898 73826 543454
rect 74382 542898 109826 543454
rect 110382 542898 145826 543454
rect 146382 542898 181826 543454
rect 182382 542898 217826 543454
rect 218382 542898 253826 543454
rect 254382 542898 289826 543454
rect 290382 542898 325826 543454
rect 326382 542898 361826 543454
rect 362382 542898 397826 543454
rect 398382 542898 433826 543454
rect 434382 542898 469826 543454
rect 470382 542898 505826 543454
rect 506382 542898 541826 543454
rect 542382 542898 577826 543454
rect 578382 542898 585342 543454
rect 585898 542898 592650 543454
rect -8726 542866 592650 542898
rect -8726 533494 592650 533526
rect -8726 532938 -8694 533494
rect -8138 532938 27866 533494
rect 28422 532938 63866 533494
rect 64422 532938 99866 533494
rect 100422 532938 135866 533494
rect 136422 532938 171866 533494
rect 172422 532938 207866 533494
rect 208422 532938 243866 533494
rect 244422 532938 279866 533494
rect 280422 532938 315866 533494
rect 316422 532938 351866 533494
rect 352422 532938 387866 533494
rect 388422 532938 423866 533494
rect 424422 532938 459866 533494
rect 460422 532938 495866 533494
rect 496422 532938 531866 533494
rect 532422 532938 567866 533494
rect 568422 532938 592062 533494
rect 592618 532938 592650 533494
rect -8726 532906 592650 532938
rect -8726 529774 592650 529806
rect -8726 529218 -7734 529774
rect -7178 529218 24146 529774
rect 24702 529218 60146 529774
rect 60702 529218 96146 529774
rect 96702 529218 132146 529774
rect 132702 529218 168146 529774
rect 168702 529218 204146 529774
rect 204702 529218 240146 529774
rect 240702 529218 276146 529774
rect 276702 529218 312146 529774
rect 312702 529218 348146 529774
rect 348702 529218 384146 529774
rect 384702 529218 420146 529774
rect 420702 529218 456146 529774
rect 456702 529218 492146 529774
rect 492702 529218 528146 529774
rect 528702 529218 564146 529774
rect 564702 529218 591102 529774
rect 591658 529218 592650 529774
rect -8726 529186 592650 529218
rect -8726 526054 592650 526086
rect -8726 525498 -6774 526054
rect -6218 525498 20426 526054
rect 20982 525498 56426 526054
rect 56982 525498 92426 526054
rect 92982 525498 128426 526054
rect 128982 525498 164426 526054
rect 164982 525498 200426 526054
rect 200982 525498 236426 526054
rect 236982 525498 272426 526054
rect 272982 525498 308426 526054
rect 308982 525498 344426 526054
rect 344982 525498 380426 526054
rect 380982 525498 416426 526054
rect 416982 525498 452426 526054
rect 452982 525498 488426 526054
rect 488982 525498 524426 526054
rect 524982 525498 560426 526054
rect 560982 525498 590142 526054
rect 590698 525498 592650 526054
rect -8726 525466 592650 525498
rect -8726 522334 592650 522366
rect -8726 521778 -5814 522334
rect -5258 521778 16706 522334
rect 17262 521778 52706 522334
rect 53262 521778 88706 522334
rect 89262 521778 124706 522334
rect 125262 521778 160706 522334
rect 161262 521778 196706 522334
rect 197262 521778 232706 522334
rect 233262 521778 268706 522334
rect 269262 521778 304706 522334
rect 305262 521778 340706 522334
rect 341262 521778 376706 522334
rect 377262 521778 412706 522334
rect 413262 521778 448706 522334
rect 449262 521778 484706 522334
rect 485262 521778 520706 522334
rect 521262 521778 556706 522334
rect 557262 521778 589182 522334
rect 589738 521778 592650 522334
rect -8726 521746 592650 521778
rect -8726 518614 592650 518646
rect -8726 518058 -4854 518614
rect -4298 518058 12986 518614
rect 13542 518058 48986 518614
rect 49542 518058 84986 518614
rect 85542 518058 120986 518614
rect 121542 518058 156986 518614
rect 157542 518058 192986 518614
rect 193542 518058 228986 518614
rect 229542 518058 264986 518614
rect 265542 518058 300986 518614
rect 301542 518058 336986 518614
rect 337542 518058 372986 518614
rect 373542 518058 408986 518614
rect 409542 518058 444986 518614
rect 445542 518058 480986 518614
rect 481542 518058 516986 518614
rect 517542 518058 552986 518614
rect 553542 518058 588222 518614
rect 588778 518058 592650 518614
rect -8726 518026 592650 518058
rect -8726 514894 592650 514926
rect -8726 514338 -3894 514894
rect -3338 514338 9266 514894
rect 9822 514338 45266 514894
rect 45822 514338 81266 514894
rect 81822 514338 117266 514894
rect 117822 514338 153266 514894
rect 153822 514338 189266 514894
rect 189822 514338 225266 514894
rect 225822 514338 261266 514894
rect 261822 514338 297266 514894
rect 297822 514338 333266 514894
rect 333822 514338 369266 514894
rect 369822 514338 405266 514894
rect 405822 514338 441266 514894
rect 441822 514338 477266 514894
rect 477822 514338 513266 514894
rect 513822 514338 549266 514894
rect 549822 514338 587262 514894
rect 587818 514338 592650 514894
rect -8726 514306 592650 514338
rect -8726 511174 592650 511206
rect -8726 510618 -2934 511174
rect -2378 510618 5546 511174
rect 6102 510618 41546 511174
rect 42102 510618 77546 511174
rect 78102 510618 113546 511174
rect 114102 510618 149546 511174
rect 150102 510618 185546 511174
rect 186102 510618 221546 511174
rect 222102 510618 257546 511174
rect 258102 510618 293546 511174
rect 294102 510618 329546 511174
rect 330102 510618 365546 511174
rect 366102 510618 401546 511174
rect 402102 510618 437546 511174
rect 438102 510618 473546 511174
rect 474102 510618 509546 511174
rect 510102 510618 545546 511174
rect 546102 510618 581546 511174
rect 582102 510618 586302 511174
rect 586858 510618 592650 511174
rect -8726 510586 592650 510618
rect -8726 507454 592650 507486
rect -8726 506898 -1974 507454
rect -1418 506898 1826 507454
rect 2382 506898 37826 507454
rect 38382 506898 73826 507454
rect 74382 506898 109826 507454
rect 110382 506898 145826 507454
rect 146382 506898 181826 507454
rect 182382 506898 217826 507454
rect 218382 506898 253826 507454
rect 254382 506898 289826 507454
rect 290382 506898 325826 507454
rect 326382 506898 361826 507454
rect 362382 506898 397826 507454
rect 398382 506898 433826 507454
rect 434382 506898 469826 507454
rect 470382 506898 505826 507454
rect 506382 506898 541826 507454
rect 542382 506898 577826 507454
rect 578382 506898 585342 507454
rect 585898 506898 592650 507454
rect -8726 506866 592650 506898
rect -8726 497494 592650 497526
rect -8726 496938 -8694 497494
rect -8138 496938 27866 497494
rect 28422 496938 63866 497494
rect 64422 496938 99866 497494
rect 100422 496938 135866 497494
rect 136422 496938 171866 497494
rect 172422 496938 207866 497494
rect 208422 496938 243866 497494
rect 244422 496938 279866 497494
rect 280422 496938 315866 497494
rect 316422 496938 351866 497494
rect 352422 496938 387866 497494
rect 388422 496938 423866 497494
rect 424422 496938 459866 497494
rect 460422 496938 495866 497494
rect 496422 496938 531866 497494
rect 532422 496938 567866 497494
rect 568422 496938 592062 497494
rect 592618 496938 592650 497494
rect -8726 496906 592650 496938
rect -8726 493774 592650 493806
rect -8726 493218 -7734 493774
rect -7178 493218 24146 493774
rect 24702 493218 60146 493774
rect 60702 493218 96146 493774
rect 96702 493218 132146 493774
rect 132702 493218 168146 493774
rect 168702 493218 204146 493774
rect 204702 493218 240146 493774
rect 240702 493218 276146 493774
rect 276702 493218 312146 493774
rect 312702 493218 348146 493774
rect 348702 493218 384146 493774
rect 384702 493218 420146 493774
rect 420702 493218 456146 493774
rect 456702 493218 492146 493774
rect 492702 493218 528146 493774
rect 528702 493218 564146 493774
rect 564702 493218 591102 493774
rect 591658 493218 592650 493774
rect -8726 493186 592650 493218
rect -8726 490054 592650 490086
rect -8726 489498 -6774 490054
rect -6218 489498 20426 490054
rect 20982 489498 56426 490054
rect 56982 489498 92426 490054
rect 92982 489498 128426 490054
rect 128982 489498 164426 490054
rect 164982 489498 200426 490054
rect 200982 489498 236426 490054
rect 236982 489498 272426 490054
rect 272982 489498 308426 490054
rect 308982 489498 344426 490054
rect 344982 489498 380426 490054
rect 380982 489498 416426 490054
rect 416982 489498 452426 490054
rect 452982 489498 488426 490054
rect 488982 489498 524426 490054
rect 524982 489498 560426 490054
rect 560982 489498 590142 490054
rect 590698 489498 592650 490054
rect -8726 489466 592650 489498
rect -8726 486334 592650 486366
rect -8726 485778 -5814 486334
rect -5258 485778 16706 486334
rect 17262 485778 52706 486334
rect 53262 485778 88706 486334
rect 89262 485778 124706 486334
rect 125262 485778 160706 486334
rect 161262 485778 196706 486334
rect 197262 485778 232706 486334
rect 233262 485778 268706 486334
rect 269262 485778 304706 486334
rect 305262 485778 340706 486334
rect 341262 485778 376706 486334
rect 377262 485778 412706 486334
rect 413262 485778 448706 486334
rect 449262 485778 484706 486334
rect 485262 485778 520706 486334
rect 521262 485778 556706 486334
rect 557262 485778 589182 486334
rect 589738 485778 592650 486334
rect -8726 485746 592650 485778
rect -8726 482614 592650 482646
rect -8726 482058 -4854 482614
rect -4298 482058 12986 482614
rect 13542 482058 48986 482614
rect 49542 482058 84986 482614
rect 85542 482058 120986 482614
rect 121542 482058 156986 482614
rect 157542 482058 192986 482614
rect 193542 482058 228986 482614
rect 229542 482058 264986 482614
rect 265542 482058 300986 482614
rect 301542 482058 336986 482614
rect 337542 482058 372986 482614
rect 373542 482058 408986 482614
rect 409542 482058 444986 482614
rect 445542 482058 480986 482614
rect 481542 482058 516986 482614
rect 517542 482058 552986 482614
rect 553542 482058 588222 482614
rect 588778 482058 592650 482614
rect -8726 482026 592650 482058
rect -8726 478894 592650 478926
rect -8726 478338 -3894 478894
rect -3338 478338 9266 478894
rect 9822 478338 45266 478894
rect 45822 478338 81266 478894
rect 81822 478338 117266 478894
rect 117822 478338 153266 478894
rect 153822 478338 189266 478894
rect 189822 478338 225266 478894
rect 225822 478338 261266 478894
rect 261822 478338 297266 478894
rect 297822 478338 333266 478894
rect 333822 478338 369266 478894
rect 369822 478338 405266 478894
rect 405822 478338 441266 478894
rect 441822 478338 477266 478894
rect 477822 478338 513266 478894
rect 513822 478338 549266 478894
rect 549822 478338 587262 478894
rect 587818 478338 592650 478894
rect -8726 478306 592650 478338
rect -8726 475174 592650 475206
rect -8726 474618 -2934 475174
rect -2378 474618 5546 475174
rect 6102 474618 41546 475174
rect 42102 474618 77546 475174
rect 78102 474618 113546 475174
rect 114102 474618 149546 475174
rect 150102 474618 185546 475174
rect 186102 474618 221546 475174
rect 222102 474618 257546 475174
rect 258102 474618 293546 475174
rect 294102 474618 329546 475174
rect 330102 474618 365546 475174
rect 366102 474618 401546 475174
rect 402102 474618 437546 475174
rect 438102 474618 473546 475174
rect 474102 474618 509546 475174
rect 510102 474618 545546 475174
rect 546102 474618 581546 475174
rect 582102 474618 586302 475174
rect 586858 474618 592650 475174
rect -8726 474586 592650 474618
rect -8726 471454 592650 471486
rect -8726 470898 -1974 471454
rect -1418 470898 1826 471454
rect 2382 470898 37826 471454
rect 38382 470898 73826 471454
rect 74382 470898 109826 471454
rect 110382 470898 145826 471454
rect 146382 470898 181826 471454
rect 182382 470898 217826 471454
rect 218382 470898 253826 471454
rect 254382 470898 289826 471454
rect 290382 470898 325826 471454
rect 326382 470898 361826 471454
rect 362382 470898 397826 471454
rect 398382 470898 433826 471454
rect 434382 470898 469826 471454
rect 470382 470898 505826 471454
rect 506382 470898 541826 471454
rect 542382 470898 577826 471454
rect 578382 470898 585342 471454
rect 585898 470898 592650 471454
rect -8726 470866 592650 470898
rect -8726 461494 592650 461526
rect -8726 460938 -8694 461494
rect -8138 460938 27866 461494
rect 28422 460938 63866 461494
rect 64422 460938 99866 461494
rect 100422 460938 135866 461494
rect 136422 460938 171866 461494
rect 172422 460938 207866 461494
rect 208422 460938 243866 461494
rect 244422 460938 279866 461494
rect 280422 460938 315866 461494
rect 316422 460938 351866 461494
rect 352422 460938 387866 461494
rect 388422 460938 423866 461494
rect 424422 460938 459866 461494
rect 460422 460938 495866 461494
rect 496422 460938 531866 461494
rect 532422 460938 567866 461494
rect 568422 460938 592062 461494
rect 592618 460938 592650 461494
rect -8726 460906 592650 460938
rect -8726 457774 592650 457806
rect -8726 457218 -7734 457774
rect -7178 457218 24146 457774
rect 24702 457218 60146 457774
rect 60702 457218 96146 457774
rect 96702 457218 132146 457774
rect 132702 457218 168146 457774
rect 168702 457218 204146 457774
rect 204702 457218 240146 457774
rect 240702 457218 276146 457774
rect 276702 457218 312146 457774
rect 312702 457218 348146 457774
rect 348702 457218 384146 457774
rect 384702 457218 420146 457774
rect 420702 457218 456146 457774
rect 456702 457218 492146 457774
rect 492702 457218 528146 457774
rect 528702 457218 564146 457774
rect 564702 457218 591102 457774
rect 591658 457218 592650 457774
rect -8726 457186 592650 457218
rect -8726 454054 592650 454086
rect -8726 453498 -6774 454054
rect -6218 453498 20426 454054
rect 20982 453498 56426 454054
rect 56982 453498 92426 454054
rect 92982 453498 128426 454054
rect 128982 453498 164426 454054
rect 164982 453498 200426 454054
rect 200982 453498 236426 454054
rect 236982 453498 272426 454054
rect 272982 453498 308426 454054
rect 308982 453498 344426 454054
rect 344982 453498 380426 454054
rect 380982 453498 416426 454054
rect 416982 453498 452426 454054
rect 452982 453498 488426 454054
rect 488982 453498 524426 454054
rect 524982 453498 560426 454054
rect 560982 453498 590142 454054
rect 590698 453498 592650 454054
rect -8726 453466 592650 453498
rect -8726 450334 592650 450366
rect -8726 449778 -5814 450334
rect -5258 449778 16706 450334
rect 17262 449778 52706 450334
rect 53262 449778 88706 450334
rect 89262 449778 124706 450334
rect 125262 449778 160706 450334
rect 161262 449778 196706 450334
rect 197262 449778 232706 450334
rect 233262 449778 268706 450334
rect 269262 449778 304706 450334
rect 305262 449778 340706 450334
rect 341262 449778 376706 450334
rect 377262 449778 412706 450334
rect 413262 449778 448706 450334
rect 449262 449778 484706 450334
rect 485262 449778 520706 450334
rect 521262 449778 556706 450334
rect 557262 449778 589182 450334
rect 589738 449778 592650 450334
rect -8726 449746 592650 449778
rect -8726 446614 592650 446646
rect -8726 446058 -4854 446614
rect -4298 446058 12986 446614
rect 13542 446058 48986 446614
rect 49542 446058 84986 446614
rect 85542 446058 120986 446614
rect 121542 446058 156986 446614
rect 157542 446058 192986 446614
rect 193542 446058 228986 446614
rect 229542 446058 264986 446614
rect 265542 446058 300986 446614
rect 301542 446058 336986 446614
rect 337542 446058 372986 446614
rect 373542 446058 408986 446614
rect 409542 446058 444986 446614
rect 445542 446058 480986 446614
rect 481542 446058 516986 446614
rect 517542 446058 552986 446614
rect 553542 446058 588222 446614
rect 588778 446058 592650 446614
rect -8726 446026 592650 446058
rect -8726 442894 592650 442926
rect -8726 442338 -3894 442894
rect -3338 442338 9266 442894
rect 9822 442338 45266 442894
rect 45822 442338 81266 442894
rect 81822 442338 117266 442894
rect 117822 442338 153266 442894
rect 153822 442338 189266 442894
rect 189822 442338 225266 442894
rect 225822 442338 261266 442894
rect 261822 442338 297266 442894
rect 297822 442338 333266 442894
rect 333822 442338 369266 442894
rect 369822 442338 405266 442894
rect 405822 442338 441266 442894
rect 441822 442338 477266 442894
rect 477822 442338 513266 442894
rect 513822 442338 549266 442894
rect 549822 442338 587262 442894
rect 587818 442338 592650 442894
rect -8726 442306 592650 442338
rect -8726 439174 592650 439206
rect -8726 438618 -2934 439174
rect -2378 438618 5546 439174
rect 6102 438618 41546 439174
rect 42102 438618 77546 439174
rect 78102 438618 113546 439174
rect 114102 438618 149546 439174
rect 150102 438618 185546 439174
rect 186102 438618 221546 439174
rect 222102 438618 257546 439174
rect 258102 438618 293546 439174
rect 294102 438618 329546 439174
rect 330102 438618 365546 439174
rect 366102 438618 401546 439174
rect 402102 438618 437546 439174
rect 438102 438618 473546 439174
rect 474102 438618 509546 439174
rect 510102 438618 545546 439174
rect 546102 438618 581546 439174
rect 582102 438618 586302 439174
rect 586858 438618 592650 439174
rect -8726 438586 592650 438618
rect -8726 435454 592650 435486
rect -8726 434898 -1974 435454
rect -1418 434898 1826 435454
rect 2382 434898 37826 435454
rect 38382 434898 73826 435454
rect 74382 434898 109826 435454
rect 110382 434898 145826 435454
rect 146382 434898 181826 435454
rect 182382 434898 217826 435454
rect 218382 434898 253826 435454
rect 254382 434898 289826 435454
rect 290382 434898 325826 435454
rect 326382 434898 361826 435454
rect 362382 434898 397826 435454
rect 398382 434898 433826 435454
rect 434382 434898 469826 435454
rect 470382 434898 505826 435454
rect 506382 434898 541826 435454
rect 542382 434898 577826 435454
rect 578382 434898 585342 435454
rect 585898 434898 592650 435454
rect -8726 434866 592650 434898
rect -8726 425494 592650 425526
rect -8726 424938 -8694 425494
rect -8138 424938 27866 425494
rect 28422 424938 63866 425494
rect 64422 424938 99866 425494
rect 100422 424938 135866 425494
rect 136422 424938 171866 425494
rect 172422 424938 207866 425494
rect 208422 424938 243866 425494
rect 244422 424938 279866 425494
rect 280422 424938 315866 425494
rect 316422 424938 351866 425494
rect 352422 424938 387866 425494
rect 388422 424938 423866 425494
rect 424422 424938 459866 425494
rect 460422 424938 495866 425494
rect 496422 424938 531866 425494
rect 532422 424938 567866 425494
rect 568422 424938 592062 425494
rect 592618 424938 592650 425494
rect -8726 424906 592650 424938
rect -8726 421774 592650 421806
rect -8726 421218 -7734 421774
rect -7178 421218 24146 421774
rect 24702 421218 60146 421774
rect 60702 421218 96146 421774
rect 96702 421218 132146 421774
rect 132702 421218 168146 421774
rect 168702 421218 204146 421774
rect 204702 421218 240146 421774
rect 240702 421218 276146 421774
rect 276702 421218 312146 421774
rect 312702 421218 348146 421774
rect 348702 421218 384146 421774
rect 384702 421218 420146 421774
rect 420702 421218 456146 421774
rect 456702 421218 492146 421774
rect 492702 421218 528146 421774
rect 528702 421218 564146 421774
rect 564702 421218 591102 421774
rect 591658 421218 592650 421774
rect -8726 421186 592650 421218
rect -8726 418054 592650 418086
rect -8726 417498 -6774 418054
rect -6218 417498 20426 418054
rect 20982 417498 56426 418054
rect 56982 417498 92426 418054
rect 92982 417498 128426 418054
rect 128982 417498 164426 418054
rect 164982 417498 200426 418054
rect 200982 417498 236426 418054
rect 236982 417498 272426 418054
rect 272982 417498 308426 418054
rect 308982 417498 344426 418054
rect 344982 417498 380426 418054
rect 380982 417498 416426 418054
rect 416982 417498 452426 418054
rect 452982 417498 488426 418054
rect 488982 417498 524426 418054
rect 524982 417498 560426 418054
rect 560982 417498 590142 418054
rect 590698 417498 592650 418054
rect -8726 417466 592650 417498
rect -8726 414334 592650 414366
rect -8726 413778 -5814 414334
rect -5258 413778 16706 414334
rect 17262 413778 52706 414334
rect 53262 413778 88706 414334
rect 89262 413778 124706 414334
rect 125262 413778 160706 414334
rect 161262 413778 196706 414334
rect 197262 413778 232706 414334
rect 233262 413778 268706 414334
rect 269262 413778 304706 414334
rect 305262 413778 340706 414334
rect 341262 413778 376706 414334
rect 377262 413778 412706 414334
rect 413262 413778 448706 414334
rect 449262 413778 484706 414334
rect 485262 413778 520706 414334
rect 521262 413778 556706 414334
rect 557262 413778 589182 414334
rect 589738 413778 592650 414334
rect -8726 413746 592650 413778
rect -8726 410614 592650 410646
rect -8726 410058 -4854 410614
rect -4298 410058 12986 410614
rect 13542 410058 48986 410614
rect 49542 410058 84986 410614
rect 85542 410058 120986 410614
rect 121542 410058 156986 410614
rect 157542 410058 192986 410614
rect 193542 410058 228986 410614
rect 229542 410058 264986 410614
rect 265542 410058 300986 410614
rect 301542 410058 336986 410614
rect 337542 410058 372986 410614
rect 373542 410058 408986 410614
rect 409542 410058 444986 410614
rect 445542 410058 480986 410614
rect 481542 410058 516986 410614
rect 517542 410058 552986 410614
rect 553542 410058 588222 410614
rect 588778 410058 592650 410614
rect -8726 410026 592650 410058
rect -8726 406894 592650 406926
rect -8726 406338 -3894 406894
rect -3338 406338 9266 406894
rect 9822 406338 45266 406894
rect 45822 406338 81266 406894
rect 81822 406338 117266 406894
rect 117822 406338 153266 406894
rect 153822 406338 189266 406894
rect 189822 406338 225266 406894
rect 225822 406338 261266 406894
rect 261822 406338 297266 406894
rect 297822 406338 333266 406894
rect 333822 406338 369266 406894
rect 369822 406338 405266 406894
rect 405822 406338 441266 406894
rect 441822 406338 477266 406894
rect 477822 406338 513266 406894
rect 513822 406338 549266 406894
rect 549822 406338 587262 406894
rect 587818 406338 592650 406894
rect -8726 406306 592650 406338
rect -8726 403174 592650 403206
rect -8726 402618 -2934 403174
rect -2378 402618 5546 403174
rect 6102 402618 41546 403174
rect 42102 402618 77546 403174
rect 78102 402618 113546 403174
rect 114102 402618 149546 403174
rect 150102 402618 185546 403174
rect 186102 402618 221546 403174
rect 222102 402618 257546 403174
rect 258102 402618 293546 403174
rect 294102 402618 329546 403174
rect 330102 402618 365546 403174
rect 366102 402618 401546 403174
rect 402102 402618 437546 403174
rect 438102 402618 473546 403174
rect 474102 402618 509546 403174
rect 510102 402618 545546 403174
rect 546102 402618 581546 403174
rect 582102 402618 586302 403174
rect 586858 402618 592650 403174
rect -8726 402586 592650 402618
rect -8726 399454 592650 399486
rect -8726 398898 -1974 399454
rect -1418 398898 1826 399454
rect 2382 398898 37826 399454
rect 38382 398898 73826 399454
rect 74382 398898 109826 399454
rect 110382 398898 145826 399454
rect 146382 398898 181826 399454
rect 182382 398898 217826 399454
rect 218382 398898 253826 399454
rect 254382 398898 289826 399454
rect 290382 398898 325826 399454
rect 326382 398898 361826 399454
rect 362382 398898 397826 399454
rect 398382 398898 433826 399454
rect 434382 398898 469826 399454
rect 470382 398898 505826 399454
rect 506382 398898 541826 399454
rect 542382 398898 577826 399454
rect 578382 398898 585342 399454
rect 585898 398898 592650 399454
rect -8726 398866 592650 398898
rect -8726 389494 592650 389526
rect -8726 388938 -8694 389494
rect -8138 388938 27866 389494
rect 28422 388938 63866 389494
rect 64422 388938 99866 389494
rect 100422 388938 135866 389494
rect 136422 388938 171866 389494
rect 172422 388938 207866 389494
rect 208422 388938 243866 389494
rect 244422 388938 279866 389494
rect 280422 388938 315866 389494
rect 316422 388938 351866 389494
rect 352422 388938 387866 389494
rect 388422 388938 423866 389494
rect 424422 388938 459866 389494
rect 460422 388938 495866 389494
rect 496422 388938 531866 389494
rect 532422 388938 567866 389494
rect 568422 388938 592062 389494
rect 592618 388938 592650 389494
rect -8726 388906 592650 388938
rect -8726 385774 592650 385806
rect -8726 385218 -7734 385774
rect -7178 385218 24146 385774
rect 24702 385218 60146 385774
rect 60702 385218 96146 385774
rect 96702 385218 132146 385774
rect 132702 385218 168146 385774
rect 168702 385218 204146 385774
rect 204702 385218 240146 385774
rect 240702 385218 276146 385774
rect 276702 385218 312146 385774
rect 312702 385218 348146 385774
rect 348702 385218 384146 385774
rect 384702 385218 420146 385774
rect 420702 385218 456146 385774
rect 456702 385218 492146 385774
rect 492702 385218 528146 385774
rect 528702 385218 564146 385774
rect 564702 385218 591102 385774
rect 591658 385218 592650 385774
rect -8726 385186 592650 385218
rect -8726 382054 592650 382086
rect -8726 381498 -6774 382054
rect -6218 381498 20426 382054
rect 20982 381498 56426 382054
rect 56982 381498 92426 382054
rect 92982 381498 128426 382054
rect 128982 381498 164426 382054
rect 164982 381498 200426 382054
rect 200982 381498 236426 382054
rect 236982 381498 272426 382054
rect 272982 381498 308426 382054
rect 308982 381498 344426 382054
rect 344982 381498 380426 382054
rect 380982 381498 416426 382054
rect 416982 381498 452426 382054
rect 452982 381498 488426 382054
rect 488982 381498 524426 382054
rect 524982 381498 560426 382054
rect 560982 381498 590142 382054
rect 590698 381498 592650 382054
rect -8726 381466 592650 381498
rect -8726 378334 592650 378366
rect -8726 377778 -5814 378334
rect -5258 377778 16706 378334
rect 17262 377778 52706 378334
rect 53262 377778 88706 378334
rect 89262 377778 124706 378334
rect 125262 377778 160706 378334
rect 161262 377778 196706 378334
rect 197262 377778 232706 378334
rect 233262 377778 268706 378334
rect 269262 377778 304706 378334
rect 305262 377778 340706 378334
rect 341262 377778 376706 378334
rect 377262 377778 412706 378334
rect 413262 377778 448706 378334
rect 449262 377778 484706 378334
rect 485262 377778 520706 378334
rect 521262 377778 556706 378334
rect 557262 377778 589182 378334
rect 589738 377778 592650 378334
rect -8726 377746 592650 377778
rect -8726 374614 592650 374646
rect -8726 374058 -4854 374614
rect -4298 374058 12986 374614
rect 13542 374058 48986 374614
rect 49542 374058 84986 374614
rect 85542 374058 120986 374614
rect 121542 374058 156986 374614
rect 157542 374058 192986 374614
rect 193542 374058 228986 374614
rect 229542 374058 264986 374614
rect 265542 374058 300986 374614
rect 301542 374058 336986 374614
rect 337542 374058 372986 374614
rect 373542 374058 408986 374614
rect 409542 374058 444986 374614
rect 445542 374058 480986 374614
rect 481542 374058 516986 374614
rect 517542 374058 552986 374614
rect 553542 374058 588222 374614
rect 588778 374058 592650 374614
rect -8726 374026 592650 374058
rect -8726 370894 592650 370926
rect -8726 370338 -3894 370894
rect -3338 370338 9266 370894
rect 9822 370338 45266 370894
rect 45822 370338 81266 370894
rect 81822 370338 117266 370894
rect 117822 370338 153266 370894
rect 153822 370338 189266 370894
rect 189822 370338 225266 370894
rect 225822 370338 261266 370894
rect 261822 370338 297266 370894
rect 297822 370338 333266 370894
rect 333822 370338 369266 370894
rect 369822 370338 405266 370894
rect 405822 370338 441266 370894
rect 441822 370338 477266 370894
rect 477822 370338 513266 370894
rect 513822 370338 549266 370894
rect 549822 370338 587262 370894
rect 587818 370338 592650 370894
rect -8726 370306 592650 370338
rect -8726 367174 592650 367206
rect -8726 366618 -2934 367174
rect -2378 366618 5546 367174
rect 6102 366618 41546 367174
rect 42102 366618 77546 367174
rect 78102 366618 113546 367174
rect 114102 366618 149546 367174
rect 150102 366618 185546 367174
rect 186102 366618 221546 367174
rect 222102 366618 257546 367174
rect 258102 366618 293546 367174
rect 294102 366618 329546 367174
rect 330102 366618 365546 367174
rect 366102 366618 401546 367174
rect 402102 366618 437546 367174
rect 438102 366618 473546 367174
rect 474102 366618 509546 367174
rect 510102 366618 545546 367174
rect 546102 366618 581546 367174
rect 582102 366618 586302 367174
rect 586858 366618 592650 367174
rect -8726 366586 592650 366618
rect -8726 363454 592650 363486
rect -8726 362898 -1974 363454
rect -1418 362898 1826 363454
rect 2382 362898 37826 363454
rect 38382 362898 73826 363454
rect 74382 362898 109826 363454
rect 110382 362898 145826 363454
rect 146382 362898 181826 363454
rect 182382 362898 217826 363454
rect 218382 362898 253826 363454
rect 254382 362898 289826 363454
rect 290382 362898 325826 363454
rect 326382 362898 361826 363454
rect 362382 362898 397826 363454
rect 398382 362898 433826 363454
rect 434382 362898 469826 363454
rect 470382 362898 505826 363454
rect 506382 362898 541826 363454
rect 542382 362898 577826 363454
rect 578382 362898 585342 363454
rect 585898 362898 592650 363454
rect -8726 362866 592650 362898
rect -8726 353494 592650 353526
rect -8726 352938 -8694 353494
rect -8138 352938 27866 353494
rect 28422 352938 63866 353494
rect 64422 352938 99866 353494
rect 100422 352938 135866 353494
rect 136422 352938 171866 353494
rect 172422 352938 207866 353494
rect 208422 352938 243866 353494
rect 244422 352938 279866 353494
rect 280422 352938 315866 353494
rect 316422 352938 351866 353494
rect 352422 352938 387866 353494
rect 388422 352938 423866 353494
rect 424422 352938 459866 353494
rect 460422 352938 495866 353494
rect 496422 352938 531866 353494
rect 532422 352938 567866 353494
rect 568422 352938 592062 353494
rect 592618 352938 592650 353494
rect -8726 352906 592650 352938
rect -8726 349774 592650 349806
rect -8726 349218 -7734 349774
rect -7178 349218 24146 349774
rect 24702 349218 60146 349774
rect 60702 349218 96146 349774
rect 96702 349218 132146 349774
rect 132702 349218 168146 349774
rect 168702 349218 204146 349774
rect 204702 349218 240146 349774
rect 240702 349218 276146 349774
rect 276702 349218 312146 349774
rect 312702 349218 348146 349774
rect 348702 349218 384146 349774
rect 384702 349218 420146 349774
rect 420702 349218 456146 349774
rect 456702 349218 492146 349774
rect 492702 349218 528146 349774
rect 528702 349218 564146 349774
rect 564702 349218 591102 349774
rect 591658 349218 592650 349774
rect -8726 349186 592650 349218
rect -8726 346054 592650 346086
rect -8726 345498 -6774 346054
rect -6218 345498 20426 346054
rect 20982 345498 56426 346054
rect 56982 345498 92426 346054
rect 92982 345498 128426 346054
rect 128982 345498 164426 346054
rect 164982 345498 200426 346054
rect 200982 345498 236426 346054
rect 236982 345498 272426 346054
rect 272982 345498 308426 346054
rect 308982 345498 344426 346054
rect 344982 345498 380426 346054
rect 380982 345498 416426 346054
rect 416982 345498 452426 346054
rect 452982 345498 488426 346054
rect 488982 345498 524426 346054
rect 524982 345498 560426 346054
rect 560982 345498 590142 346054
rect 590698 345498 592650 346054
rect -8726 345466 592650 345498
rect -8726 342334 592650 342366
rect -8726 341778 -5814 342334
rect -5258 341778 16706 342334
rect 17262 341778 52706 342334
rect 53262 341778 88706 342334
rect 89262 341778 124706 342334
rect 125262 341778 160706 342334
rect 161262 341778 196706 342334
rect 197262 341778 232706 342334
rect 233262 341778 268706 342334
rect 269262 341778 304706 342334
rect 305262 341778 340706 342334
rect 341262 341778 376706 342334
rect 377262 341778 412706 342334
rect 413262 341778 448706 342334
rect 449262 341778 484706 342334
rect 485262 341778 520706 342334
rect 521262 341778 556706 342334
rect 557262 341778 589182 342334
rect 589738 341778 592650 342334
rect -8726 341746 592650 341778
rect -8726 338614 592650 338646
rect -8726 338058 -4854 338614
rect -4298 338058 12986 338614
rect 13542 338058 48986 338614
rect 49542 338058 84986 338614
rect 85542 338058 120986 338614
rect 121542 338058 156986 338614
rect 157542 338058 192986 338614
rect 193542 338058 228986 338614
rect 229542 338058 264986 338614
rect 265542 338058 300986 338614
rect 301542 338058 336986 338614
rect 337542 338058 372986 338614
rect 373542 338058 408986 338614
rect 409542 338058 444986 338614
rect 445542 338058 480986 338614
rect 481542 338058 516986 338614
rect 517542 338058 552986 338614
rect 553542 338058 588222 338614
rect 588778 338058 592650 338614
rect -8726 338026 592650 338058
rect -8726 334894 592650 334926
rect -8726 334338 -3894 334894
rect -3338 334338 9266 334894
rect 9822 334338 45266 334894
rect 45822 334338 81266 334894
rect 81822 334338 117266 334894
rect 117822 334338 153266 334894
rect 153822 334338 189266 334894
rect 189822 334338 225266 334894
rect 225822 334338 261266 334894
rect 261822 334338 297266 334894
rect 297822 334338 333266 334894
rect 333822 334338 369266 334894
rect 369822 334338 405266 334894
rect 405822 334338 441266 334894
rect 441822 334338 477266 334894
rect 477822 334338 513266 334894
rect 513822 334338 549266 334894
rect 549822 334338 587262 334894
rect 587818 334338 592650 334894
rect -8726 334306 592650 334338
rect -8726 331174 592650 331206
rect -8726 330618 -2934 331174
rect -2378 330618 5546 331174
rect 6102 330618 41546 331174
rect 42102 330618 77546 331174
rect 78102 330618 113546 331174
rect 114102 330618 149546 331174
rect 150102 330618 185546 331174
rect 186102 330618 221546 331174
rect 222102 330618 257546 331174
rect 258102 330618 293546 331174
rect 294102 330618 329546 331174
rect 330102 330618 365546 331174
rect 366102 330618 401546 331174
rect 402102 330618 437546 331174
rect 438102 330618 473546 331174
rect 474102 330618 509546 331174
rect 510102 330618 545546 331174
rect 546102 330618 581546 331174
rect 582102 330618 586302 331174
rect 586858 330618 592650 331174
rect -8726 330586 592650 330618
rect -8726 327454 592650 327486
rect -8726 326898 -1974 327454
rect -1418 326898 1826 327454
rect 2382 326898 37826 327454
rect 38382 326898 73826 327454
rect 74382 326898 109826 327454
rect 110382 326898 145826 327454
rect 146382 326898 181826 327454
rect 182382 326898 217826 327454
rect 218382 326898 253826 327454
rect 254382 326898 289826 327454
rect 290382 326898 325826 327454
rect 326382 326898 361826 327454
rect 362382 326898 397826 327454
rect 398382 326898 433826 327454
rect 434382 326898 469826 327454
rect 470382 326898 505826 327454
rect 506382 326898 541826 327454
rect 542382 326898 577826 327454
rect 578382 326898 585342 327454
rect 585898 326898 592650 327454
rect -8726 326866 592650 326898
rect -8726 317494 592650 317526
rect -8726 316938 -8694 317494
rect -8138 316938 27866 317494
rect 28422 316938 63866 317494
rect 64422 316938 99866 317494
rect 100422 316938 135866 317494
rect 136422 316938 171866 317494
rect 172422 316938 207866 317494
rect 208422 316938 243866 317494
rect 244422 316938 279866 317494
rect 280422 316938 315866 317494
rect 316422 316938 351866 317494
rect 352422 316938 387866 317494
rect 388422 316938 423866 317494
rect 424422 316938 459866 317494
rect 460422 316938 495866 317494
rect 496422 316938 531866 317494
rect 532422 316938 567866 317494
rect 568422 316938 592062 317494
rect 592618 316938 592650 317494
rect -8726 316906 592650 316938
rect -8726 313774 592650 313806
rect -8726 313218 -7734 313774
rect -7178 313218 24146 313774
rect 24702 313218 60146 313774
rect 60702 313218 96146 313774
rect 96702 313218 132146 313774
rect 132702 313218 168146 313774
rect 168702 313218 204146 313774
rect 204702 313218 240146 313774
rect 240702 313218 276146 313774
rect 276702 313218 312146 313774
rect 312702 313218 348146 313774
rect 348702 313218 384146 313774
rect 384702 313218 420146 313774
rect 420702 313218 456146 313774
rect 456702 313218 492146 313774
rect 492702 313218 528146 313774
rect 528702 313218 564146 313774
rect 564702 313218 591102 313774
rect 591658 313218 592650 313774
rect -8726 313186 592650 313218
rect -8726 310054 592650 310086
rect -8726 309498 -6774 310054
rect -6218 309498 20426 310054
rect 20982 309498 56426 310054
rect 56982 309498 92426 310054
rect 92982 309498 128426 310054
rect 128982 309498 164426 310054
rect 164982 309498 200426 310054
rect 200982 309498 236426 310054
rect 236982 309498 272426 310054
rect 272982 309498 308426 310054
rect 308982 309498 344426 310054
rect 344982 309498 380426 310054
rect 380982 309498 416426 310054
rect 416982 309498 452426 310054
rect 452982 309498 488426 310054
rect 488982 309498 524426 310054
rect 524982 309498 560426 310054
rect 560982 309498 590142 310054
rect 590698 309498 592650 310054
rect -8726 309466 592650 309498
rect -8726 306334 592650 306366
rect -8726 305778 -5814 306334
rect -5258 305778 16706 306334
rect 17262 305778 52706 306334
rect 53262 305778 88706 306334
rect 89262 305778 124706 306334
rect 125262 305778 160706 306334
rect 161262 305778 196706 306334
rect 197262 305778 232706 306334
rect 233262 305778 268706 306334
rect 269262 305778 304706 306334
rect 305262 305778 340706 306334
rect 341262 305778 376706 306334
rect 377262 305778 412706 306334
rect 413262 305778 448706 306334
rect 449262 305778 484706 306334
rect 485262 305778 520706 306334
rect 521262 305778 556706 306334
rect 557262 305778 589182 306334
rect 589738 305778 592650 306334
rect -8726 305746 592650 305778
rect -8726 302614 592650 302646
rect -8726 302058 -4854 302614
rect -4298 302058 12986 302614
rect 13542 302058 48986 302614
rect 49542 302058 84986 302614
rect 85542 302058 120986 302614
rect 121542 302058 156986 302614
rect 157542 302058 192986 302614
rect 193542 302058 228986 302614
rect 229542 302058 264986 302614
rect 265542 302058 300986 302614
rect 301542 302058 336986 302614
rect 337542 302058 372986 302614
rect 373542 302058 408986 302614
rect 409542 302058 444986 302614
rect 445542 302058 480986 302614
rect 481542 302058 516986 302614
rect 517542 302058 552986 302614
rect 553542 302058 588222 302614
rect 588778 302058 592650 302614
rect -8726 302026 592650 302058
rect -8726 298894 592650 298926
rect -8726 298338 -3894 298894
rect -3338 298338 9266 298894
rect 9822 298338 45266 298894
rect 45822 298338 81266 298894
rect 81822 298338 117266 298894
rect 117822 298338 153266 298894
rect 153822 298338 189266 298894
rect 189822 298338 225266 298894
rect 225822 298338 261266 298894
rect 261822 298338 297266 298894
rect 297822 298338 333266 298894
rect 333822 298338 369266 298894
rect 369822 298338 405266 298894
rect 405822 298338 441266 298894
rect 441822 298338 477266 298894
rect 477822 298338 513266 298894
rect 513822 298338 549266 298894
rect 549822 298338 587262 298894
rect 587818 298338 592650 298894
rect -8726 298306 592650 298338
rect -8726 295174 592650 295206
rect -8726 294618 -2934 295174
rect -2378 294618 5546 295174
rect 6102 294618 41546 295174
rect 42102 294618 77546 295174
rect 78102 294618 113546 295174
rect 114102 294618 149546 295174
rect 150102 294618 185546 295174
rect 186102 294618 221546 295174
rect 222102 294618 257546 295174
rect 258102 294618 293546 295174
rect 294102 294618 329546 295174
rect 330102 294618 365546 295174
rect 366102 294618 401546 295174
rect 402102 294618 437546 295174
rect 438102 294618 473546 295174
rect 474102 294618 509546 295174
rect 510102 294618 545546 295174
rect 546102 294618 581546 295174
rect 582102 294618 586302 295174
rect 586858 294618 592650 295174
rect -8726 294586 592650 294618
rect -8726 291454 592650 291486
rect -8726 290898 -1974 291454
rect -1418 290898 1826 291454
rect 2382 290898 37826 291454
rect 38382 290898 73826 291454
rect 74382 290898 109826 291454
rect 110382 290898 145826 291454
rect 146382 290898 181826 291454
rect 182382 290898 217826 291454
rect 218382 290898 253826 291454
rect 254382 290898 289826 291454
rect 290382 290898 325826 291454
rect 326382 290898 361826 291454
rect 362382 290898 397826 291454
rect 398382 290898 433826 291454
rect 434382 290898 469826 291454
rect 470382 290898 505826 291454
rect 506382 290898 541826 291454
rect 542382 290898 577826 291454
rect 578382 290898 585342 291454
rect 585898 290898 592650 291454
rect -8726 290866 592650 290898
rect -8726 281494 592650 281526
rect -8726 280938 -8694 281494
rect -8138 280938 27866 281494
rect 28422 280938 63866 281494
rect 64422 280938 99866 281494
rect 100422 280938 135866 281494
rect 136422 280938 171866 281494
rect 172422 280938 243866 281494
rect 244422 280938 279866 281494
rect 280422 280938 315866 281494
rect 316422 280938 351866 281494
rect 352422 280938 387866 281494
rect 388422 280938 423866 281494
rect 424422 280938 459866 281494
rect 460422 280938 495866 281494
rect 496422 280938 531866 281494
rect 532422 280938 567866 281494
rect 568422 280938 592062 281494
rect 592618 280938 592650 281494
rect -8726 280906 592650 280938
rect -8726 277774 592650 277806
rect -8726 277218 -7734 277774
rect -7178 277218 60146 277774
rect 60702 277218 96146 277774
rect 96702 277218 132146 277774
rect 132702 277218 168146 277774
rect 168702 277218 204146 277774
rect 204702 277218 240146 277774
rect 240702 277218 276146 277774
rect 276702 277218 312146 277774
rect 312702 277218 348146 277774
rect 348702 277218 384146 277774
rect 384702 277218 420146 277774
rect 420702 277218 456146 277774
rect 456702 277218 492146 277774
rect 492702 277218 528146 277774
rect 528702 277218 564146 277774
rect 564702 277218 591102 277774
rect 591658 277218 592650 277774
rect -8726 277186 592650 277218
rect -8726 274054 592650 274086
rect -8726 273498 -6774 274054
rect -6218 273498 20426 274054
rect 20982 273818 39290 274054
rect 39526 273818 56426 274054
rect 20982 273734 56426 273818
rect 20982 273498 39290 273734
rect 39526 273498 56426 273734
rect 56982 273818 70010 274054
rect 70246 273818 100730 274054
rect 100966 273818 128426 274054
rect 56982 273734 128426 273818
rect 56982 273498 70010 273734
rect 70246 273498 100730 273734
rect 100966 273498 128426 273734
rect 128982 273818 131450 274054
rect 131686 273818 162170 274054
rect 162406 273818 164426 274054
rect 128982 273734 164426 273818
rect 128982 273498 131450 273734
rect 131686 273498 162170 273734
rect 162406 273498 164426 273734
rect 164982 273818 192890 274054
rect 193126 273818 223610 274054
rect 223846 273818 236426 274054
rect 164982 273734 236426 273818
rect 164982 273498 192890 273734
rect 193126 273498 223610 273734
rect 223846 273498 236426 273734
rect 236982 273818 254330 274054
rect 254566 273818 272426 274054
rect 236982 273734 272426 273818
rect 236982 273498 254330 273734
rect 254566 273498 272426 273734
rect 272982 273818 285050 274054
rect 285286 273818 308426 274054
rect 272982 273734 308426 273818
rect 272982 273498 285050 273734
rect 285286 273498 308426 273734
rect 308982 273498 344426 274054
rect 344982 273498 380426 274054
rect 380982 273498 416426 274054
rect 416982 273498 452426 274054
rect 452982 273498 488426 274054
rect 488982 273498 524426 274054
rect 524982 273498 560426 274054
rect 560982 273498 590142 274054
rect 590698 273498 592650 274054
rect -8726 273466 592650 273498
rect -8726 270334 592650 270366
rect -8726 269778 -5814 270334
rect -5258 269778 16706 270334
rect 17262 270098 31610 270334
rect 31846 270098 52706 270334
rect 17262 270014 52706 270098
rect 17262 269778 31610 270014
rect 31846 269778 52706 270014
rect 53262 270098 62330 270334
rect 62566 270098 88706 270334
rect 53262 270014 88706 270098
rect 53262 269778 62330 270014
rect 62566 269778 88706 270014
rect 89262 270098 93050 270334
rect 93286 270098 123770 270334
rect 124006 270098 124706 270334
rect 89262 270014 124706 270098
rect 89262 269778 93050 270014
rect 93286 269778 123770 270014
rect 124006 269778 124706 270014
rect 125262 270098 154490 270334
rect 154726 270098 160706 270334
rect 125262 270014 160706 270098
rect 125262 269778 154490 270014
rect 154726 269778 160706 270014
rect 161262 270098 185210 270334
rect 185446 270098 196706 270334
rect 161262 270014 196706 270098
rect 161262 269778 185210 270014
rect 185446 269778 196706 270014
rect 197262 270098 215930 270334
rect 216166 270098 232706 270334
rect 197262 270014 232706 270098
rect 197262 269778 215930 270014
rect 216166 269778 232706 270014
rect 233262 270098 246650 270334
rect 246886 270098 268706 270334
rect 233262 270014 268706 270098
rect 233262 269778 246650 270014
rect 246886 269778 268706 270014
rect 269262 270098 277370 270334
rect 277606 270098 304706 270334
rect 269262 270014 304706 270098
rect 269262 269778 277370 270014
rect 277606 269778 304706 270014
rect 305262 269778 340706 270334
rect 341262 269778 376706 270334
rect 377262 269778 412706 270334
rect 413262 269778 448706 270334
rect 449262 269778 484706 270334
rect 485262 269778 520706 270334
rect 521262 269778 556706 270334
rect 557262 269778 589182 270334
rect 589738 269778 592650 270334
rect -8726 269746 592650 269778
rect -8726 266614 592650 266646
rect -8726 266058 -4854 266614
rect -4298 266058 12986 266614
rect 13542 266058 48986 266614
rect 49542 266058 120986 266614
rect 121542 266058 156986 266614
rect 157542 266058 228986 266614
rect 229542 266058 264986 266614
rect 265542 266058 300986 266614
rect 301542 266058 336986 266614
rect 337542 266058 372986 266614
rect 373542 266058 408986 266614
rect 409542 266058 444986 266614
rect 445542 266058 480986 266614
rect 481542 266058 516986 266614
rect 517542 266058 552986 266614
rect 553542 266058 588222 266614
rect 588778 266058 592650 266614
rect -8726 266026 592650 266058
rect -8726 262894 592650 262926
rect -8726 262338 -3894 262894
rect -3338 262338 9266 262894
rect 9822 262338 45266 262894
rect 45822 262338 81266 262894
rect 81822 262338 117266 262894
rect 117822 262338 153266 262894
rect 153822 262338 189266 262894
rect 189822 262338 225266 262894
rect 225822 262338 297266 262894
rect 297822 262338 333266 262894
rect 333822 262338 369266 262894
rect 369822 262338 405266 262894
rect 405822 262338 441266 262894
rect 441822 262338 477266 262894
rect 477822 262338 513266 262894
rect 513822 262338 549266 262894
rect 549822 262338 587262 262894
rect 587818 262338 592650 262894
rect -8726 262306 592650 262338
rect -8726 259174 592650 259206
rect -8726 258618 -2934 259174
rect -2378 258618 5546 259174
rect 6102 258938 23930 259174
rect 24166 258938 41546 259174
rect 6102 258854 41546 258938
rect 6102 258618 23930 258854
rect 24166 258618 41546 258854
rect 42102 258938 54650 259174
rect 54886 258938 85370 259174
rect 85606 258938 113546 259174
rect 42102 258854 113546 258938
rect 42102 258618 54650 258854
rect 54886 258618 85370 258854
rect 85606 258618 113546 258854
rect 114102 258938 116090 259174
rect 116326 258938 146810 259174
rect 147046 258938 149546 259174
rect 114102 258854 149546 258938
rect 114102 258618 116090 258854
rect 116326 258618 146810 258854
rect 147046 258618 149546 258854
rect 150102 258938 177530 259174
rect 177766 258938 208250 259174
rect 208486 258938 221546 259174
rect 150102 258854 221546 258938
rect 150102 258618 177530 258854
rect 177766 258618 208250 258854
rect 208486 258618 221546 258854
rect 222102 258938 238970 259174
rect 239206 258938 257546 259174
rect 222102 258854 257546 258938
rect 222102 258618 238970 258854
rect 239206 258618 257546 258854
rect 258102 258938 269690 259174
rect 269926 258938 293546 259174
rect 258102 258854 293546 258938
rect 258102 258618 269690 258854
rect 269926 258618 293546 258854
rect 294102 258618 329546 259174
rect 330102 258618 365546 259174
rect 366102 258618 401546 259174
rect 402102 258618 437546 259174
rect 438102 258618 473546 259174
rect 474102 258618 509546 259174
rect 510102 258618 545546 259174
rect 546102 258618 581546 259174
rect 582102 258618 586302 259174
rect 586858 258618 592650 259174
rect -8726 258586 592650 258618
rect -8726 255454 592650 255486
rect -8726 254898 -1974 255454
rect -1418 254898 1826 255454
rect 2382 255218 16250 255454
rect 16486 255218 37826 255454
rect 2382 255134 37826 255218
rect 2382 254898 16250 255134
rect 16486 254898 37826 255134
rect 38382 255218 46970 255454
rect 47206 255218 73826 255454
rect 38382 255134 73826 255218
rect 38382 254898 46970 255134
rect 47206 254898 73826 255134
rect 74382 255218 77690 255454
rect 77926 255218 108410 255454
rect 108646 255218 109826 255454
rect 74382 255134 109826 255218
rect 74382 254898 77690 255134
rect 77926 254898 108410 255134
rect 108646 254898 109826 255134
rect 110382 255218 139130 255454
rect 139366 255218 145826 255454
rect 110382 255134 145826 255218
rect 110382 254898 139130 255134
rect 139366 254898 145826 255134
rect 146382 255218 169850 255454
rect 170086 255218 181826 255454
rect 146382 255134 181826 255218
rect 146382 254898 169850 255134
rect 170086 254898 181826 255134
rect 182382 255218 200570 255454
rect 200806 255218 217826 255454
rect 182382 255134 217826 255218
rect 182382 254898 200570 255134
rect 200806 254898 217826 255134
rect 218382 255218 231290 255454
rect 231526 255218 262010 255454
rect 262246 255218 289826 255454
rect 218382 255134 289826 255218
rect 218382 254898 231290 255134
rect 231526 254898 262010 255134
rect 262246 254898 289826 255134
rect 290382 254898 325826 255454
rect 326382 254898 361826 255454
rect 362382 254898 397826 255454
rect 398382 254898 433826 255454
rect 434382 254898 469826 255454
rect 470382 254898 505826 255454
rect 506382 254898 541826 255454
rect 542382 254898 577826 255454
rect 578382 254898 585342 255454
rect 585898 254898 592650 255454
rect -8726 254866 592650 254898
rect -8726 245494 592650 245526
rect -8726 244938 -8694 245494
rect -8138 244938 27866 245494
rect 28422 244938 63866 245494
rect 64422 244938 99866 245494
rect 100422 244938 135866 245494
rect 136422 244938 171866 245494
rect 172422 244938 243866 245494
rect 244422 244938 279866 245494
rect 280422 244938 315866 245494
rect 316422 244938 351866 245494
rect 352422 244938 387866 245494
rect 388422 244938 423866 245494
rect 424422 244938 459866 245494
rect 460422 244938 495866 245494
rect 496422 244938 531866 245494
rect 532422 244938 567866 245494
rect 568422 244938 592062 245494
rect 592618 244938 592650 245494
rect -8726 244906 592650 244938
rect -8726 241774 592650 241806
rect -8726 241218 -7734 241774
rect -7178 241218 60146 241774
rect 60702 241218 96146 241774
rect 96702 241218 132146 241774
rect 132702 241218 168146 241774
rect 168702 241218 204146 241774
rect 204702 241218 240146 241774
rect 240702 241218 276146 241774
rect 276702 241218 312146 241774
rect 312702 241218 348146 241774
rect 348702 241218 384146 241774
rect 384702 241218 420146 241774
rect 420702 241218 456146 241774
rect 456702 241218 492146 241774
rect 492702 241218 528146 241774
rect 528702 241218 564146 241774
rect 564702 241218 591102 241774
rect 591658 241218 592650 241774
rect -8726 241186 592650 241218
rect -8726 238054 592650 238086
rect -8726 237498 -6774 238054
rect -6218 237498 20426 238054
rect 20982 237818 39290 238054
rect 39526 237818 56426 238054
rect 20982 237734 56426 237818
rect 20982 237498 39290 237734
rect 39526 237498 56426 237734
rect 56982 237818 70010 238054
rect 70246 237818 100730 238054
rect 100966 237818 128426 238054
rect 56982 237734 128426 237818
rect 56982 237498 70010 237734
rect 70246 237498 100730 237734
rect 100966 237498 128426 237734
rect 128982 237818 131450 238054
rect 131686 237818 162170 238054
rect 162406 237818 164426 238054
rect 128982 237734 164426 237818
rect 128982 237498 131450 237734
rect 131686 237498 162170 237734
rect 162406 237498 164426 237734
rect 164982 237818 192890 238054
rect 193126 237818 223610 238054
rect 223846 237818 236426 238054
rect 164982 237734 236426 237818
rect 164982 237498 192890 237734
rect 193126 237498 223610 237734
rect 223846 237498 236426 237734
rect 236982 237818 254330 238054
rect 254566 237818 272426 238054
rect 236982 237734 272426 237818
rect 236982 237498 254330 237734
rect 254566 237498 272426 237734
rect 272982 237818 285050 238054
rect 285286 237818 308426 238054
rect 272982 237734 308426 237818
rect 272982 237498 285050 237734
rect 285286 237498 308426 237734
rect 308982 237498 344426 238054
rect 344982 237498 380426 238054
rect 380982 237498 416426 238054
rect 416982 237498 452426 238054
rect 452982 237498 488426 238054
rect 488982 237498 524426 238054
rect 524982 237498 560426 238054
rect 560982 237498 590142 238054
rect 590698 237498 592650 238054
rect -8726 237466 592650 237498
rect -8726 234334 592650 234366
rect -8726 233778 -5814 234334
rect -5258 233778 16706 234334
rect 17262 234098 31610 234334
rect 31846 234098 52706 234334
rect 17262 234014 52706 234098
rect 17262 233778 31610 234014
rect 31846 233778 52706 234014
rect 53262 234098 62330 234334
rect 62566 234098 88706 234334
rect 53262 234014 88706 234098
rect 53262 233778 62330 234014
rect 62566 233778 88706 234014
rect 89262 234098 93050 234334
rect 93286 234098 123770 234334
rect 124006 234098 124706 234334
rect 89262 234014 124706 234098
rect 89262 233778 93050 234014
rect 93286 233778 123770 234014
rect 124006 233778 124706 234014
rect 125262 234098 154490 234334
rect 154726 234098 160706 234334
rect 125262 234014 160706 234098
rect 125262 233778 154490 234014
rect 154726 233778 160706 234014
rect 161262 234098 185210 234334
rect 185446 234098 196706 234334
rect 161262 234014 196706 234098
rect 161262 233778 185210 234014
rect 185446 233778 196706 234014
rect 197262 234098 215930 234334
rect 216166 234098 232706 234334
rect 197262 234014 232706 234098
rect 197262 233778 215930 234014
rect 216166 233778 232706 234014
rect 233262 234098 246650 234334
rect 246886 234098 268706 234334
rect 233262 234014 268706 234098
rect 233262 233778 246650 234014
rect 246886 233778 268706 234014
rect 269262 234098 277370 234334
rect 277606 234098 304706 234334
rect 269262 234014 304706 234098
rect 269262 233778 277370 234014
rect 277606 233778 304706 234014
rect 305262 233778 340706 234334
rect 341262 233778 376706 234334
rect 377262 233778 412706 234334
rect 413262 233778 448706 234334
rect 449262 233778 484706 234334
rect 485262 233778 520706 234334
rect 521262 233778 556706 234334
rect 557262 233778 589182 234334
rect 589738 233778 592650 234334
rect -8726 233746 592650 233778
rect -8726 230614 592650 230646
rect -8726 230058 -4854 230614
rect -4298 230058 12986 230614
rect 13542 230058 48986 230614
rect 49542 230058 120986 230614
rect 121542 230058 156986 230614
rect 157542 230058 228986 230614
rect 229542 230058 264986 230614
rect 265542 230058 300986 230614
rect 301542 230058 336986 230614
rect 337542 230058 372986 230614
rect 373542 230058 408986 230614
rect 409542 230058 444986 230614
rect 445542 230058 480986 230614
rect 481542 230058 516986 230614
rect 517542 230058 552986 230614
rect 553542 230058 588222 230614
rect 588778 230058 592650 230614
rect -8726 230026 592650 230058
rect -8726 226894 592650 226926
rect -8726 226338 -3894 226894
rect -3338 226338 9266 226894
rect 9822 226338 45266 226894
rect 45822 226338 81266 226894
rect 81822 226338 117266 226894
rect 117822 226338 153266 226894
rect 153822 226338 189266 226894
rect 189822 226338 225266 226894
rect 225822 226338 297266 226894
rect 297822 226338 333266 226894
rect 333822 226338 369266 226894
rect 369822 226338 405266 226894
rect 405822 226338 441266 226894
rect 441822 226338 477266 226894
rect 477822 226338 513266 226894
rect 513822 226338 549266 226894
rect 549822 226338 587262 226894
rect 587818 226338 592650 226894
rect -8726 226306 592650 226338
rect -8726 223174 592650 223206
rect -8726 222618 -2934 223174
rect -2378 222618 5546 223174
rect 6102 222938 23930 223174
rect 24166 222938 41546 223174
rect 6102 222854 41546 222938
rect 6102 222618 23930 222854
rect 24166 222618 41546 222854
rect 42102 222938 54650 223174
rect 54886 222938 85370 223174
rect 85606 222938 113546 223174
rect 42102 222854 113546 222938
rect 42102 222618 54650 222854
rect 54886 222618 85370 222854
rect 85606 222618 113546 222854
rect 114102 222938 116090 223174
rect 116326 222938 146810 223174
rect 147046 222938 149546 223174
rect 114102 222854 149546 222938
rect 114102 222618 116090 222854
rect 116326 222618 146810 222854
rect 147046 222618 149546 222854
rect 150102 222938 177530 223174
rect 177766 222938 208250 223174
rect 208486 222938 221546 223174
rect 150102 222854 221546 222938
rect 150102 222618 177530 222854
rect 177766 222618 208250 222854
rect 208486 222618 221546 222854
rect 222102 222938 238970 223174
rect 239206 222938 257546 223174
rect 222102 222854 257546 222938
rect 222102 222618 238970 222854
rect 239206 222618 257546 222854
rect 258102 222938 269690 223174
rect 269926 222938 293546 223174
rect 258102 222854 293546 222938
rect 258102 222618 269690 222854
rect 269926 222618 293546 222854
rect 294102 222618 329546 223174
rect 330102 222618 365546 223174
rect 366102 222618 401546 223174
rect 402102 222618 437546 223174
rect 438102 222618 473546 223174
rect 474102 222618 509546 223174
rect 510102 222618 545546 223174
rect 546102 222618 581546 223174
rect 582102 222618 586302 223174
rect 586858 222618 592650 223174
rect -8726 222586 592650 222618
rect -8726 219454 592650 219486
rect -8726 218898 -1974 219454
rect -1418 218898 1826 219454
rect 2382 219218 16250 219454
rect 16486 219218 37826 219454
rect 2382 219134 37826 219218
rect 2382 218898 16250 219134
rect 16486 218898 37826 219134
rect 38382 219218 46970 219454
rect 47206 219218 73826 219454
rect 38382 219134 73826 219218
rect 38382 218898 46970 219134
rect 47206 218898 73826 219134
rect 74382 219218 77690 219454
rect 77926 219218 108410 219454
rect 108646 219218 109826 219454
rect 74382 219134 109826 219218
rect 74382 218898 77690 219134
rect 77926 218898 108410 219134
rect 108646 218898 109826 219134
rect 110382 219218 139130 219454
rect 139366 219218 145826 219454
rect 110382 219134 145826 219218
rect 110382 218898 139130 219134
rect 139366 218898 145826 219134
rect 146382 219218 169850 219454
rect 170086 219218 181826 219454
rect 146382 219134 181826 219218
rect 146382 218898 169850 219134
rect 170086 218898 181826 219134
rect 182382 219218 200570 219454
rect 200806 219218 217826 219454
rect 182382 219134 217826 219218
rect 182382 218898 200570 219134
rect 200806 218898 217826 219134
rect 218382 219218 231290 219454
rect 231526 219218 262010 219454
rect 262246 219218 289826 219454
rect 218382 219134 289826 219218
rect 218382 218898 231290 219134
rect 231526 218898 262010 219134
rect 262246 218898 289826 219134
rect 290382 218898 325826 219454
rect 326382 218898 361826 219454
rect 362382 218898 397826 219454
rect 398382 218898 433826 219454
rect 434382 218898 469826 219454
rect 470382 218898 505826 219454
rect 506382 218898 541826 219454
rect 542382 218898 577826 219454
rect 578382 218898 585342 219454
rect 585898 218898 592650 219454
rect -8726 218866 592650 218898
rect -8726 209494 592650 209526
rect -8726 208938 -8694 209494
rect -8138 208938 27866 209494
rect 28422 208938 63866 209494
rect 64422 208938 99866 209494
rect 100422 208938 135866 209494
rect 136422 208938 171866 209494
rect 172422 208938 243866 209494
rect 244422 208938 279866 209494
rect 280422 208938 315866 209494
rect 316422 208938 351866 209494
rect 352422 208938 387866 209494
rect 388422 208938 423866 209494
rect 424422 208938 459866 209494
rect 460422 208938 495866 209494
rect 496422 208938 531866 209494
rect 532422 208938 567866 209494
rect 568422 208938 592062 209494
rect 592618 208938 592650 209494
rect -8726 208906 592650 208938
rect -8726 205774 592650 205806
rect -8726 205218 -7734 205774
rect -7178 205218 60146 205774
rect 60702 205218 96146 205774
rect 96702 205218 132146 205774
rect 132702 205218 168146 205774
rect 168702 205218 204146 205774
rect 204702 205218 240146 205774
rect 240702 205218 276146 205774
rect 276702 205218 312146 205774
rect 312702 205218 348146 205774
rect 348702 205218 384146 205774
rect 384702 205218 420146 205774
rect 420702 205218 456146 205774
rect 456702 205218 492146 205774
rect 492702 205218 528146 205774
rect 528702 205218 564146 205774
rect 564702 205218 591102 205774
rect 591658 205218 592650 205774
rect -8726 205186 592650 205218
rect -8726 202054 592650 202086
rect -8726 201498 -6774 202054
rect -6218 201498 20426 202054
rect 20982 201818 39290 202054
rect 39526 201818 56426 202054
rect 20982 201734 56426 201818
rect 20982 201498 39290 201734
rect 39526 201498 56426 201734
rect 56982 201818 70010 202054
rect 70246 201818 100730 202054
rect 100966 201818 128426 202054
rect 56982 201734 128426 201818
rect 56982 201498 70010 201734
rect 70246 201498 100730 201734
rect 100966 201498 128426 201734
rect 128982 201818 131450 202054
rect 131686 201818 162170 202054
rect 162406 201818 164426 202054
rect 128982 201734 164426 201818
rect 128982 201498 131450 201734
rect 131686 201498 162170 201734
rect 162406 201498 164426 201734
rect 164982 201818 192890 202054
rect 193126 201818 223610 202054
rect 223846 201818 236426 202054
rect 164982 201734 236426 201818
rect 164982 201498 192890 201734
rect 193126 201498 223610 201734
rect 223846 201498 236426 201734
rect 236982 201818 254330 202054
rect 254566 201818 272426 202054
rect 236982 201734 272426 201818
rect 236982 201498 254330 201734
rect 254566 201498 272426 201734
rect 272982 201818 285050 202054
rect 285286 201818 308426 202054
rect 272982 201734 308426 201818
rect 272982 201498 285050 201734
rect 285286 201498 308426 201734
rect 308982 201498 344426 202054
rect 344982 201498 380426 202054
rect 380982 201498 416426 202054
rect 416982 201498 452426 202054
rect 452982 201498 488426 202054
rect 488982 201498 524426 202054
rect 524982 201498 560426 202054
rect 560982 201498 590142 202054
rect 590698 201498 592650 202054
rect -8726 201466 592650 201498
rect -8726 198334 592650 198366
rect -8726 197778 -5814 198334
rect -5258 197778 16706 198334
rect 17262 198098 31610 198334
rect 31846 198098 52706 198334
rect 17262 198014 52706 198098
rect 17262 197778 31610 198014
rect 31846 197778 52706 198014
rect 53262 198098 62330 198334
rect 62566 198098 88706 198334
rect 53262 198014 88706 198098
rect 53262 197778 62330 198014
rect 62566 197778 88706 198014
rect 89262 198098 93050 198334
rect 93286 198098 123770 198334
rect 124006 198098 124706 198334
rect 89262 198014 124706 198098
rect 89262 197778 93050 198014
rect 93286 197778 123770 198014
rect 124006 197778 124706 198014
rect 125262 198098 154490 198334
rect 154726 198098 160706 198334
rect 125262 198014 160706 198098
rect 125262 197778 154490 198014
rect 154726 197778 160706 198014
rect 161262 198098 185210 198334
rect 185446 198098 196706 198334
rect 161262 198014 196706 198098
rect 161262 197778 185210 198014
rect 185446 197778 196706 198014
rect 197262 198098 215930 198334
rect 216166 198098 232706 198334
rect 197262 198014 232706 198098
rect 197262 197778 215930 198014
rect 216166 197778 232706 198014
rect 233262 198098 246650 198334
rect 246886 198098 268706 198334
rect 233262 198014 268706 198098
rect 233262 197778 246650 198014
rect 246886 197778 268706 198014
rect 269262 198098 277370 198334
rect 277606 198098 304706 198334
rect 269262 198014 304706 198098
rect 269262 197778 277370 198014
rect 277606 197778 304706 198014
rect 305262 197778 340706 198334
rect 341262 197778 376706 198334
rect 377262 197778 412706 198334
rect 413262 197778 448706 198334
rect 449262 197778 484706 198334
rect 485262 197778 520706 198334
rect 521262 197778 556706 198334
rect 557262 197778 589182 198334
rect 589738 197778 592650 198334
rect -8726 197746 592650 197778
rect -8726 194614 592650 194646
rect -8726 194058 -4854 194614
rect -4298 194058 12986 194614
rect 13542 194058 48986 194614
rect 49542 194058 120986 194614
rect 121542 194058 156986 194614
rect 157542 194058 228986 194614
rect 229542 194058 264986 194614
rect 265542 194058 300986 194614
rect 301542 194058 336986 194614
rect 337542 194058 372986 194614
rect 373542 194058 408986 194614
rect 409542 194058 444986 194614
rect 445542 194058 480986 194614
rect 481542 194058 516986 194614
rect 517542 194058 552986 194614
rect 553542 194058 588222 194614
rect 588778 194058 592650 194614
rect -8726 194026 592650 194058
rect -8726 190894 592650 190926
rect -8726 190338 -3894 190894
rect -3338 190338 9266 190894
rect 9822 190338 45266 190894
rect 45822 190338 81266 190894
rect 81822 190338 117266 190894
rect 117822 190338 153266 190894
rect 153822 190338 189266 190894
rect 189822 190338 225266 190894
rect 225822 190338 297266 190894
rect 297822 190338 333266 190894
rect 333822 190338 369266 190894
rect 369822 190338 405266 190894
rect 405822 190338 441266 190894
rect 441822 190338 477266 190894
rect 477822 190338 513266 190894
rect 513822 190338 549266 190894
rect 549822 190338 587262 190894
rect 587818 190338 592650 190894
rect -8726 190306 592650 190338
rect -8726 187174 592650 187206
rect -8726 186618 -2934 187174
rect -2378 186618 5546 187174
rect 6102 186938 23930 187174
rect 24166 186938 41546 187174
rect 6102 186854 41546 186938
rect 6102 186618 23930 186854
rect 24166 186618 41546 186854
rect 42102 186938 54650 187174
rect 54886 186938 85370 187174
rect 85606 186938 113546 187174
rect 42102 186854 113546 186938
rect 42102 186618 54650 186854
rect 54886 186618 85370 186854
rect 85606 186618 113546 186854
rect 114102 186938 116090 187174
rect 116326 186938 146810 187174
rect 147046 186938 149546 187174
rect 114102 186854 149546 186938
rect 114102 186618 116090 186854
rect 116326 186618 146810 186854
rect 147046 186618 149546 186854
rect 150102 186938 177530 187174
rect 177766 186938 208250 187174
rect 208486 186938 221546 187174
rect 150102 186854 221546 186938
rect 150102 186618 177530 186854
rect 177766 186618 208250 186854
rect 208486 186618 221546 186854
rect 222102 186938 238970 187174
rect 239206 186938 257546 187174
rect 222102 186854 257546 186938
rect 222102 186618 238970 186854
rect 239206 186618 257546 186854
rect 258102 186938 269690 187174
rect 269926 186938 293546 187174
rect 258102 186854 293546 186938
rect 258102 186618 269690 186854
rect 269926 186618 293546 186854
rect 294102 186618 329546 187174
rect 330102 186618 365546 187174
rect 366102 186618 401546 187174
rect 402102 186618 437546 187174
rect 438102 186618 473546 187174
rect 474102 186618 509546 187174
rect 510102 186618 545546 187174
rect 546102 186618 581546 187174
rect 582102 186618 586302 187174
rect 586858 186618 592650 187174
rect -8726 186586 592650 186618
rect -8726 183454 592650 183486
rect -8726 182898 -1974 183454
rect -1418 182898 1826 183454
rect 2382 183218 16250 183454
rect 16486 183218 37826 183454
rect 2382 183134 37826 183218
rect 2382 182898 16250 183134
rect 16486 182898 37826 183134
rect 38382 183218 46970 183454
rect 47206 183218 73826 183454
rect 38382 183134 73826 183218
rect 38382 182898 46970 183134
rect 47206 182898 73826 183134
rect 74382 183218 77690 183454
rect 77926 183218 108410 183454
rect 108646 183218 109826 183454
rect 74382 183134 109826 183218
rect 74382 182898 77690 183134
rect 77926 182898 108410 183134
rect 108646 182898 109826 183134
rect 110382 183218 139130 183454
rect 139366 183218 145826 183454
rect 110382 183134 145826 183218
rect 110382 182898 139130 183134
rect 139366 182898 145826 183134
rect 146382 183218 169850 183454
rect 170086 183218 181826 183454
rect 146382 183134 181826 183218
rect 146382 182898 169850 183134
rect 170086 182898 181826 183134
rect 182382 183218 200570 183454
rect 200806 183218 217826 183454
rect 182382 183134 217826 183218
rect 182382 182898 200570 183134
rect 200806 182898 217826 183134
rect 218382 183218 231290 183454
rect 231526 183218 262010 183454
rect 262246 183218 289826 183454
rect 218382 183134 289826 183218
rect 218382 182898 231290 183134
rect 231526 182898 262010 183134
rect 262246 182898 289826 183134
rect 290382 182898 325826 183454
rect 326382 182898 361826 183454
rect 362382 182898 397826 183454
rect 398382 182898 433826 183454
rect 434382 182898 469826 183454
rect 470382 182898 505826 183454
rect 506382 182898 541826 183454
rect 542382 182898 577826 183454
rect 578382 182898 585342 183454
rect 585898 182898 592650 183454
rect -8726 182866 592650 182898
rect -8726 173494 592650 173526
rect -8726 172938 -8694 173494
rect -8138 172938 27866 173494
rect 28422 172938 63866 173494
rect 64422 172938 99866 173494
rect 100422 172938 135866 173494
rect 136422 172938 171866 173494
rect 172422 172938 243866 173494
rect 244422 172938 279866 173494
rect 280422 172938 315866 173494
rect 316422 172938 351866 173494
rect 352422 172938 387866 173494
rect 388422 172938 423866 173494
rect 424422 172938 459866 173494
rect 460422 172938 495866 173494
rect 496422 172938 531866 173494
rect 532422 172938 567866 173494
rect 568422 172938 592062 173494
rect 592618 172938 592650 173494
rect -8726 172906 592650 172938
rect -8726 169774 592650 169806
rect -8726 169218 -7734 169774
rect -7178 169218 60146 169774
rect 60702 169218 96146 169774
rect 96702 169218 132146 169774
rect 132702 169218 168146 169774
rect 168702 169218 204146 169774
rect 204702 169218 240146 169774
rect 240702 169218 276146 169774
rect 276702 169218 312146 169774
rect 312702 169218 348146 169774
rect 348702 169218 384146 169774
rect 384702 169218 420146 169774
rect 420702 169218 456146 169774
rect 456702 169218 492146 169774
rect 492702 169218 528146 169774
rect 528702 169218 564146 169774
rect 564702 169218 591102 169774
rect 591658 169218 592650 169774
rect -8726 169186 592650 169218
rect -8726 166054 592650 166086
rect -8726 165498 -6774 166054
rect -6218 165498 20426 166054
rect 20982 165818 39290 166054
rect 39526 165818 56426 166054
rect 20982 165734 56426 165818
rect 20982 165498 39290 165734
rect 39526 165498 56426 165734
rect 56982 165818 70010 166054
rect 70246 165818 100730 166054
rect 100966 165818 128426 166054
rect 56982 165734 128426 165818
rect 56982 165498 70010 165734
rect 70246 165498 100730 165734
rect 100966 165498 128426 165734
rect 128982 165818 131450 166054
rect 131686 165818 162170 166054
rect 162406 165818 164426 166054
rect 128982 165734 164426 165818
rect 128982 165498 131450 165734
rect 131686 165498 162170 165734
rect 162406 165498 164426 165734
rect 164982 165818 192890 166054
rect 193126 165818 223610 166054
rect 223846 165818 236426 166054
rect 164982 165734 236426 165818
rect 164982 165498 192890 165734
rect 193126 165498 223610 165734
rect 223846 165498 236426 165734
rect 236982 165818 254330 166054
rect 254566 165818 272426 166054
rect 236982 165734 272426 165818
rect 236982 165498 254330 165734
rect 254566 165498 272426 165734
rect 272982 165818 285050 166054
rect 285286 165818 308426 166054
rect 272982 165734 308426 165818
rect 272982 165498 285050 165734
rect 285286 165498 308426 165734
rect 308982 165498 344426 166054
rect 344982 165498 380426 166054
rect 380982 165498 416426 166054
rect 416982 165498 452426 166054
rect 452982 165498 488426 166054
rect 488982 165498 524426 166054
rect 524982 165498 560426 166054
rect 560982 165498 590142 166054
rect 590698 165498 592650 166054
rect -8726 165466 592650 165498
rect -8726 162334 592650 162366
rect -8726 161778 -5814 162334
rect -5258 161778 16706 162334
rect 17262 162098 31610 162334
rect 31846 162098 52706 162334
rect 17262 162014 52706 162098
rect 17262 161778 31610 162014
rect 31846 161778 52706 162014
rect 53262 162098 62330 162334
rect 62566 162098 88706 162334
rect 53262 162014 88706 162098
rect 53262 161778 62330 162014
rect 62566 161778 88706 162014
rect 89262 162098 93050 162334
rect 93286 162098 123770 162334
rect 124006 162098 124706 162334
rect 89262 162014 124706 162098
rect 89262 161778 93050 162014
rect 93286 161778 123770 162014
rect 124006 161778 124706 162014
rect 125262 162098 154490 162334
rect 154726 162098 160706 162334
rect 125262 162014 160706 162098
rect 125262 161778 154490 162014
rect 154726 161778 160706 162014
rect 161262 162098 185210 162334
rect 185446 162098 196706 162334
rect 161262 162014 196706 162098
rect 161262 161778 185210 162014
rect 185446 161778 196706 162014
rect 197262 162098 215930 162334
rect 216166 162098 232706 162334
rect 197262 162014 232706 162098
rect 197262 161778 215930 162014
rect 216166 161778 232706 162014
rect 233262 162098 246650 162334
rect 246886 162098 268706 162334
rect 233262 162014 268706 162098
rect 233262 161778 246650 162014
rect 246886 161778 268706 162014
rect 269262 162098 277370 162334
rect 277606 162098 304706 162334
rect 269262 162014 304706 162098
rect 269262 161778 277370 162014
rect 277606 161778 304706 162014
rect 305262 161778 340706 162334
rect 341262 161778 376706 162334
rect 377262 161778 412706 162334
rect 413262 161778 448706 162334
rect 449262 161778 484706 162334
rect 485262 161778 520706 162334
rect 521262 161778 556706 162334
rect 557262 161778 589182 162334
rect 589738 161778 592650 162334
rect -8726 161746 592650 161778
rect -8726 158614 592650 158646
rect -8726 158058 -4854 158614
rect -4298 158058 12986 158614
rect 13542 158058 48986 158614
rect 49542 158058 120986 158614
rect 121542 158058 156986 158614
rect 157542 158058 228986 158614
rect 229542 158058 264986 158614
rect 265542 158058 300986 158614
rect 301542 158058 336986 158614
rect 337542 158058 372986 158614
rect 373542 158058 408986 158614
rect 409542 158058 444986 158614
rect 445542 158058 480986 158614
rect 481542 158058 516986 158614
rect 517542 158058 552986 158614
rect 553542 158058 588222 158614
rect 588778 158058 592650 158614
rect -8726 158026 592650 158058
rect -8726 154894 592650 154926
rect -8726 154338 -3894 154894
rect -3338 154338 9266 154894
rect 9822 154338 45266 154894
rect 45822 154338 81266 154894
rect 81822 154338 117266 154894
rect 117822 154338 153266 154894
rect 153822 154338 189266 154894
rect 189822 154338 225266 154894
rect 225822 154338 297266 154894
rect 297822 154338 333266 154894
rect 333822 154338 369266 154894
rect 369822 154338 405266 154894
rect 405822 154338 441266 154894
rect 441822 154338 477266 154894
rect 477822 154338 513266 154894
rect 513822 154338 549266 154894
rect 549822 154338 587262 154894
rect 587818 154338 592650 154894
rect -8726 154306 592650 154338
rect -8726 151174 592650 151206
rect -8726 150618 -2934 151174
rect -2378 150618 5546 151174
rect 6102 150938 23930 151174
rect 24166 150938 41546 151174
rect 6102 150854 41546 150938
rect 6102 150618 23930 150854
rect 24166 150618 41546 150854
rect 42102 150938 54650 151174
rect 54886 150938 85370 151174
rect 85606 150938 113546 151174
rect 42102 150854 113546 150938
rect 42102 150618 54650 150854
rect 54886 150618 85370 150854
rect 85606 150618 113546 150854
rect 114102 150938 116090 151174
rect 116326 150938 146810 151174
rect 147046 150938 149546 151174
rect 114102 150854 149546 150938
rect 114102 150618 116090 150854
rect 116326 150618 146810 150854
rect 147046 150618 149546 150854
rect 150102 150938 177530 151174
rect 177766 150938 208250 151174
rect 208486 150938 221546 151174
rect 150102 150854 221546 150938
rect 150102 150618 177530 150854
rect 177766 150618 208250 150854
rect 208486 150618 221546 150854
rect 222102 150938 238970 151174
rect 239206 150938 257546 151174
rect 222102 150854 257546 150938
rect 222102 150618 238970 150854
rect 239206 150618 257546 150854
rect 258102 150938 269690 151174
rect 269926 150938 293546 151174
rect 258102 150854 293546 150938
rect 258102 150618 269690 150854
rect 269926 150618 293546 150854
rect 294102 150618 329546 151174
rect 330102 150618 365546 151174
rect 366102 150618 401546 151174
rect 402102 150618 437546 151174
rect 438102 150618 473546 151174
rect 474102 150618 509546 151174
rect 510102 150618 545546 151174
rect 546102 150618 581546 151174
rect 582102 150618 586302 151174
rect 586858 150618 592650 151174
rect -8726 150586 592650 150618
rect -8726 147454 592650 147486
rect -8726 146898 -1974 147454
rect -1418 146898 1826 147454
rect 2382 147218 16250 147454
rect 16486 147218 37826 147454
rect 2382 147134 37826 147218
rect 2382 146898 16250 147134
rect 16486 146898 37826 147134
rect 38382 147218 46970 147454
rect 47206 147218 73826 147454
rect 38382 147134 73826 147218
rect 38382 146898 46970 147134
rect 47206 146898 73826 147134
rect 74382 147218 77690 147454
rect 77926 147218 108410 147454
rect 108646 147218 109826 147454
rect 74382 147134 109826 147218
rect 74382 146898 77690 147134
rect 77926 146898 108410 147134
rect 108646 146898 109826 147134
rect 110382 147218 139130 147454
rect 139366 147218 145826 147454
rect 110382 147134 145826 147218
rect 110382 146898 139130 147134
rect 139366 146898 145826 147134
rect 146382 147218 169850 147454
rect 170086 147218 181826 147454
rect 146382 147134 181826 147218
rect 146382 146898 169850 147134
rect 170086 146898 181826 147134
rect 182382 147218 200570 147454
rect 200806 147218 217826 147454
rect 182382 147134 217826 147218
rect 182382 146898 200570 147134
rect 200806 146898 217826 147134
rect 218382 147218 231290 147454
rect 231526 147218 262010 147454
rect 262246 147218 289826 147454
rect 218382 147134 289826 147218
rect 218382 146898 231290 147134
rect 231526 146898 262010 147134
rect 262246 146898 289826 147134
rect 290382 146898 325826 147454
rect 326382 146898 361826 147454
rect 362382 146898 397826 147454
rect 398382 146898 433826 147454
rect 434382 146898 469826 147454
rect 470382 146898 505826 147454
rect 506382 146898 541826 147454
rect 542382 146898 577826 147454
rect 578382 146898 585342 147454
rect 585898 146898 592650 147454
rect -8726 146866 592650 146898
rect -8726 137494 592650 137526
rect -8726 136938 -8694 137494
rect -8138 136938 27866 137494
rect 28422 136938 63866 137494
rect 64422 136938 99866 137494
rect 100422 136938 135866 137494
rect 136422 136938 171866 137494
rect 172422 136938 243866 137494
rect 244422 136938 279866 137494
rect 280422 136938 315866 137494
rect 316422 136938 351866 137494
rect 352422 136938 387866 137494
rect 388422 136938 423866 137494
rect 424422 136938 459866 137494
rect 460422 136938 495866 137494
rect 496422 136938 531866 137494
rect 532422 136938 567866 137494
rect 568422 136938 592062 137494
rect 592618 136938 592650 137494
rect -8726 136906 592650 136938
rect -8726 133774 592650 133806
rect -8726 133218 -7734 133774
rect -7178 133218 60146 133774
rect 60702 133218 96146 133774
rect 96702 133218 132146 133774
rect 132702 133218 168146 133774
rect 168702 133218 204146 133774
rect 204702 133218 240146 133774
rect 240702 133218 276146 133774
rect 276702 133218 312146 133774
rect 312702 133218 348146 133774
rect 348702 133218 384146 133774
rect 384702 133218 420146 133774
rect 420702 133218 456146 133774
rect 456702 133218 492146 133774
rect 492702 133218 528146 133774
rect 528702 133218 564146 133774
rect 564702 133218 591102 133774
rect 591658 133218 592650 133774
rect -8726 133186 592650 133218
rect -8726 130054 592650 130086
rect -8726 129498 -6774 130054
rect -6218 129498 20426 130054
rect 20982 129818 39290 130054
rect 39526 129818 56426 130054
rect 20982 129734 56426 129818
rect 20982 129498 39290 129734
rect 39526 129498 56426 129734
rect 56982 129818 70010 130054
rect 70246 129818 100730 130054
rect 100966 129818 128426 130054
rect 56982 129734 128426 129818
rect 56982 129498 70010 129734
rect 70246 129498 100730 129734
rect 100966 129498 128426 129734
rect 128982 129818 131450 130054
rect 131686 129818 162170 130054
rect 162406 129818 164426 130054
rect 128982 129734 164426 129818
rect 128982 129498 131450 129734
rect 131686 129498 162170 129734
rect 162406 129498 164426 129734
rect 164982 129818 192890 130054
rect 193126 129818 223610 130054
rect 223846 129818 236426 130054
rect 164982 129734 236426 129818
rect 164982 129498 192890 129734
rect 193126 129498 223610 129734
rect 223846 129498 236426 129734
rect 236982 129818 254330 130054
rect 254566 129818 272426 130054
rect 236982 129734 272426 129818
rect 236982 129498 254330 129734
rect 254566 129498 272426 129734
rect 272982 129818 285050 130054
rect 285286 129818 308426 130054
rect 272982 129734 308426 129818
rect 272982 129498 285050 129734
rect 285286 129498 308426 129734
rect 308982 129498 344426 130054
rect 344982 129498 380426 130054
rect 380982 129498 416426 130054
rect 416982 129498 452426 130054
rect 452982 129498 488426 130054
rect 488982 129498 524426 130054
rect 524982 129498 560426 130054
rect 560982 129498 590142 130054
rect 590698 129498 592650 130054
rect -8726 129466 592650 129498
rect -8726 126334 592650 126366
rect -8726 125778 -5814 126334
rect -5258 126098 31610 126334
rect 31846 126098 52706 126334
rect -5258 126014 52706 126098
rect -5258 125778 31610 126014
rect 31846 125778 52706 126014
rect 53262 126098 62330 126334
rect 62566 126098 88706 126334
rect 53262 126014 88706 126098
rect 53262 125778 62330 126014
rect 62566 125778 88706 126014
rect 89262 126098 93050 126334
rect 93286 126098 123770 126334
rect 124006 126098 124706 126334
rect 89262 126014 124706 126098
rect 89262 125778 93050 126014
rect 93286 125778 123770 126014
rect 124006 125778 124706 126014
rect 125262 126098 154490 126334
rect 154726 126098 160706 126334
rect 125262 126014 160706 126098
rect 125262 125778 154490 126014
rect 154726 125778 160706 126014
rect 161262 126098 185210 126334
rect 185446 126098 196706 126334
rect 161262 126014 196706 126098
rect 161262 125778 185210 126014
rect 185446 125778 196706 126014
rect 197262 126098 215930 126334
rect 216166 126098 232706 126334
rect 197262 126014 232706 126098
rect 197262 125778 215930 126014
rect 216166 125778 232706 126014
rect 233262 126098 246650 126334
rect 246886 126098 268706 126334
rect 233262 126014 268706 126098
rect 233262 125778 246650 126014
rect 246886 125778 268706 126014
rect 269262 126098 277370 126334
rect 277606 126098 304706 126334
rect 269262 126014 304706 126098
rect 269262 125778 277370 126014
rect 277606 125778 304706 126014
rect 305262 125778 340706 126334
rect 341262 125778 376706 126334
rect 377262 125778 412706 126334
rect 413262 125778 448706 126334
rect 449262 125778 484706 126334
rect 485262 125778 520706 126334
rect 521262 125778 556706 126334
rect 557262 125778 589182 126334
rect 589738 125778 592650 126334
rect -8726 125746 592650 125778
rect -8726 122614 592650 122646
rect -8726 122058 -4854 122614
rect -4298 122058 12986 122614
rect 13542 122058 48986 122614
rect 49542 122058 120986 122614
rect 121542 122058 156986 122614
rect 157542 122058 228986 122614
rect 229542 122058 264986 122614
rect 265542 122058 300986 122614
rect 301542 122058 336986 122614
rect 337542 122058 372986 122614
rect 373542 122058 408986 122614
rect 409542 122058 444986 122614
rect 445542 122058 480986 122614
rect 481542 122058 516986 122614
rect 517542 122058 552986 122614
rect 553542 122058 588222 122614
rect 588778 122058 592650 122614
rect -8726 122026 592650 122058
rect -8726 118894 592650 118926
rect -8726 118338 -3894 118894
rect -3338 118338 9266 118894
rect 9822 118338 45266 118894
rect 45822 118338 81266 118894
rect 81822 118338 117266 118894
rect 117822 118338 153266 118894
rect 153822 118338 189266 118894
rect 189822 118338 225266 118894
rect 225822 118338 297266 118894
rect 297822 118338 333266 118894
rect 333822 118338 369266 118894
rect 369822 118338 405266 118894
rect 405822 118338 441266 118894
rect 441822 118338 477266 118894
rect 477822 118338 513266 118894
rect 513822 118338 549266 118894
rect 549822 118338 587262 118894
rect 587818 118338 592650 118894
rect -8726 118306 592650 118338
rect -8726 115174 592650 115206
rect -8726 114618 -2934 115174
rect -2378 114618 5546 115174
rect 6102 114938 17310 115174
rect 17546 114938 23930 115174
rect 24166 114938 41546 115174
rect 6102 114854 41546 114938
rect 6102 114618 17310 114854
rect 17546 114618 23930 114854
rect 24166 114618 41546 114854
rect 42102 114938 54650 115174
rect 54886 114938 85370 115174
rect 85606 114938 116090 115174
rect 116326 114938 146810 115174
rect 147046 114938 149546 115174
rect 42102 114854 149546 114938
rect 42102 114618 54650 114854
rect 54886 114618 85370 114854
rect 85606 114618 116090 114854
rect 116326 114618 146810 114854
rect 147046 114618 149546 114854
rect 150102 114938 177530 115174
rect 177766 114938 208250 115174
rect 208486 114938 221546 115174
rect 150102 114854 221546 114938
rect 150102 114618 177530 114854
rect 177766 114618 208250 114854
rect 208486 114618 221546 114854
rect 222102 114938 238970 115174
rect 239206 114938 257546 115174
rect 222102 114854 257546 114938
rect 222102 114618 238970 114854
rect 239206 114618 257546 114854
rect 258102 114938 269690 115174
rect 269926 114938 293546 115174
rect 258102 114854 293546 114938
rect 258102 114618 269690 114854
rect 269926 114618 293546 114854
rect 294102 114618 329546 115174
rect 330102 114618 365546 115174
rect 366102 114618 401546 115174
rect 402102 114618 437546 115174
rect 438102 114618 473546 115174
rect 474102 114618 509546 115174
rect 510102 114618 545546 115174
rect 546102 114618 581546 115174
rect 582102 114618 586302 115174
rect 586858 114618 592650 115174
rect -8726 114586 592650 114618
rect -8726 111454 592650 111486
rect -8726 110898 -1974 111454
rect -1418 110898 1826 111454
rect 2382 111218 16250 111454
rect 16486 111218 37826 111454
rect 2382 111134 37826 111218
rect 2382 110898 16250 111134
rect 16486 110898 37826 111134
rect 38382 111218 46970 111454
rect 47206 111218 73826 111454
rect 38382 111134 73826 111218
rect 38382 110898 46970 111134
rect 47206 110898 73826 111134
rect 74382 111218 77690 111454
rect 77926 111218 108410 111454
rect 108646 111218 109826 111454
rect 74382 111134 109826 111218
rect 74382 110898 77690 111134
rect 77926 110898 108410 111134
rect 108646 110898 109826 111134
rect 110382 111218 139130 111454
rect 139366 111218 145826 111454
rect 110382 111134 145826 111218
rect 110382 110898 139130 111134
rect 139366 110898 145826 111134
rect 146382 111218 169850 111454
rect 170086 111218 181826 111454
rect 146382 111134 181826 111218
rect 146382 110898 169850 111134
rect 170086 110898 181826 111134
rect 182382 111218 200570 111454
rect 200806 111218 217826 111454
rect 182382 111134 217826 111218
rect 182382 110898 200570 111134
rect 200806 110898 217826 111134
rect 218382 111218 231290 111454
rect 231526 111218 262010 111454
rect 262246 111218 289826 111454
rect 218382 111134 289826 111218
rect 218382 110898 231290 111134
rect 231526 110898 262010 111134
rect 262246 110898 289826 111134
rect 290382 110898 325826 111454
rect 326382 110898 361826 111454
rect 362382 110898 397826 111454
rect 398382 110898 433826 111454
rect 434382 110898 469826 111454
rect 470382 110898 505826 111454
rect 506382 110898 541826 111454
rect 542382 110898 577826 111454
rect 578382 110898 585342 111454
rect 585898 110898 592650 111454
rect -8726 110866 592650 110898
rect -8726 101494 592650 101526
rect -8726 100938 -8694 101494
rect -8138 100938 27866 101494
rect 28422 100938 63866 101494
rect 64422 100938 99866 101494
rect 100422 100938 135866 101494
rect 136422 100938 171866 101494
rect 172422 100938 243866 101494
rect 244422 100938 279866 101494
rect 280422 100938 315866 101494
rect 316422 100938 351866 101494
rect 352422 100938 387866 101494
rect 388422 100938 423866 101494
rect 424422 100938 459866 101494
rect 460422 100938 495866 101494
rect 496422 100938 531866 101494
rect 532422 100938 567866 101494
rect 568422 100938 592062 101494
rect 592618 100938 592650 101494
rect -8726 100906 592650 100938
rect -8726 97774 592650 97806
rect -8726 97218 -7734 97774
rect -7178 97218 60146 97774
rect 60702 97218 96146 97774
rect 96702 97218 132146 97774
rect 132702 97218 168146 97774
rect 168702 97218 204146 97774
rect 204702 97218 240146 97774
rect 240702 97218 276146 97774
rect 276702 97218 312146 97774
rect 312702 97218 348146 97774
rect 348702 97218 384146 97774
rect 384702 97218 420146 97774
rect 420702 97218 456146 97774
rect 456702 97218 492146 97774
rect 492702 97218 528146 97774
rect 528702 97218 564146 97774
rect 564702 97218 591102 97774
rect 591658 97218 592650 97774
rect -8726 97186 592650 97218
rect -8726 94054 592650 94086
rect -8726 93498 -6774 94054
rect -6218 93498 20426 94054
rect 20982 93818 39290 94054
rect 39526 93818 56426 94054
rect 20982 93734 56426 93818
rect 20982 93498 39290 93734
rect 39526 93498 56426 93734
rect 56982 93818 70010 94054
rect 70246 93818 100730 94054
rect 100966 93818 128426 94054
rect 56982 93734 128426 93818
rect 56982 93498 70010 93734
rect 70246 93498 100730 93734
rect 100966 93498 128426 93734
rect 128982 93818 131450 94054
rect 131686 93818 162170 94054
rect 162406 93818 164426 94054
rect 128982 93734 164426 93818
rect 128982 93498 131450 93734
rect 131686 93498 162170 93734
rect 162406 93498 164426 93734
rect 164982 93818 192890 94054
rect 193126 93818 223610 94054
rect 223846 93818 236426 94054
rect 164982 93734 236426 93818
rect 164982 93498 192890 93734
rect 193126 93498 223610 93734
rect 223846 93498 236426 93734
rect 236982 93818 254330 94054
rect 254566 93818 272426 94054
rect 236982 93734 272426 93818
rect 236982 93498 254330 93734
rect 254566 93498 272426 93734
rect 272982 93818 285050 94054
rect 285286 93818 308426 94054
rect 272982 93734 308426 93818
rect 272982 93498 285050 93734
rect 285286 93498 308426 93734
rect 308982 93498 344426 94054
rect 344982 93498 380426 94054
rect 380982 93498 416426 94054
rect 416982 93498 452426 94054
rect 452982 93498 488426 94054
rect 488982 93498 524426 94054
rect 524982 93498 560426 94054
rect 560982 93498 590142 94054
rect 590698 93498 592650 94054
rect -8726 93466 592650 93498
rect -8726 90334 592650 90366
rect -8726 89778 -5814 90334
rect -5258 90098 31610 90334
rect 31846 90098 52706 90334
rect -5258 90014 52706 90098
rect -5258 89778 31610 90014
rect 31846 89778 52706 90014
rect 53262 90098 62330 90334
rect 62566 90098 88706 90334
rect 53262 90014 88706 90098
rect 53262 89778 62330 90014
rect 62566 89778 88706 90014
rect 89262 90098 93050 90334
rect 93286 90098 123770 90334
rect 124006 90098 124706 90334
rect 89262 90014 124706 90098
rect 89262 89778 93050 90014
rect 93286 89778 123770 90014
rect 124006 89778 124706 90014
rect 125262 90098 154490 90334
rect 154726 90098 160706 90334
rect 125262 90014 160706 90098
rect 125262 89778 154490 90014
rect 154726 89778 160706 90014
rect 161262 90098 185210 90334
rect 185446 90098 196706 90334
rect 161262 90014 196706 90098
rect 161262 89778 185210 90014
rect 185446 89778 196706 90014
rect 197262 90098 215930 90334
rect 216166 90098 232706 90334
rect 197262 90014 232706 90098
rect 197262 89778 215930 90014
rect 216166 89778 232706 90014
rect 233262 90098 246650 90334
rect 246886 90098 268706 90334
rect 233262 90014 268706 90098
rect 233262 89778 246650 90014
rect 246886 89778 268706 90014
rect 269262 90098 277370 90334
rect 277606 90098 304706 90334
rect 269262 90014 304706 90098
rect 269262 89778 277370 90014
rect 277606 89778 304706 90014
rect 305262 89778 340706 90334
rect 341262 89778 376706 90334
rect 377262 89778 412706 90334
rect 413262 89778 448706 90334
rect 449262 89778 484706 90334
rect 485262 89778 520706 90334
rect 521262 89778 556706 90334
rect 557262 89778 589182 90334
rect 589738 89778 592650 90334
rect -8726 89746 592650 89778
rect -8726 86614 592650 86646
rect -8726 86058 -4854 86614
rect -4298 86058 12986 86614
rect 13542 86058 48986 86614
rect 49542 86058 120986 86614
rect 121542 86058 156986 86614
rect 157542 86058 228986 86614
rect 229542 86058 264986 86614
rect 265542 86058 300986 86614
rect 301542 86058 336986 86614
rect 337542 86058 372986 86614
rect 373542 86058 408986 86614
rect 409542 86058 444986 86614
rect 445542 86058 480986 86614
rect 481542 86058 516986 86614
rect 517542 86058 552986 86614
rect 553542 86058 588222 86614
rect 588778 86058 592650 86614
rect -8726 86026 592650 86058
rect -8726 82894 592650 82926
rect -8726 82338 -3894 82894
rect -3338 82338 9266 82894
rect 9822 82338 45266 82894
rect 45822 82338 81266 82894
rect 81822 82338 117266 82894
rect 117822 82338 153266 82894
rect 153822 82338 189266 82894
rect 189822 82338 225266 82894
rect 225822 82338 297266 82894
rect 297822 82338 333266 82894
rect 333822 82338 369266 82894
rect 369822 82338 405266 82894
rect 405822 82338 441266 82894
rect 441822 82338 477266 82894
rect 477822 82338 513266 82894
rect 513822 82338 549266 82894
rect 549822 82338 587262 82894
rect 587818 82338 592650 82894
rect -8726 82306 592650 82338
rect -8726 79174 592650 79206
rect -8726 78618 -2934 79174
rect -2378 78618 5546 79174
rect 6102 78938 17310 79174
rect 17546 78938 23930 79174
rect 24166 78938 41546 79174
rect 6102 78854 41546 78938
rect 6102 78618 17310 78854
rect 17546 78618 23930 78854
rect 24166 78618 41546 78854
rect 42102 78938 54650 79174
rect 54886 78938 85370 79174
rect 85606 78938 116090 79174
rect 116326 78938 146810 79174
rect 147046 78938 149546 79174
rect 42102 78854 149546 78938
rect 42102 78618 54650 78854
rect 54886 78618 85370 78854
rect 85606 78618 116090 78854
rect 116326 78618 146810 78854
rect 147046 78618 149546 78854
rect 150102 78938 177530 79174
rect 177766 78938 208250 79174
rect 208486 78938 221546 79174
rect 150102 78854 221546 78938
rect 150102 78618 177530 78854
rect 177766 78618 208250 78854
rect 208486 78618 221546 78854
rect 222102 78938 238970 79174
rect 239206 78938 257546 79174
rect 222102 78854 257546 78938
rect 222102 78618 238970 78854
rect 239206 78618 257546 78854
rect 258102 78938 269690 79174
rect 269926 78938 293546 79174
rect 258102 78854 293546 78938
rect 258102 78618 269690 78854
rect 269926 78618 293546 78854
rect 294102 78618 329546 79174
rect 330102 78618 365546 79174
rect 366102 78618 401546 79174
rect 402102 78618 437546 79174
rect 438102 78618 473546 79174
rect 474102 78618 509546 79174
rect 510102 78618 545546 79174
rect 546102 78618 581546 79174
rect 582102 78618 586302 79174
rect 586858 78618 592650 79174
rect -8726 78586 592650 78618
rect -8726 75454 592650 75486
rect -8726 74898 -1974 75454
rect -1418 74898 1826 75454
rect 2382 75218 16250 75454
rect 16486 75218 37826 75454
rect 2382 75134 37826 75218
rect 2382 74898 16250 75134
rect 16486 74898 37826 75134
rect 38382 75218 46970 75454
rect 47206 75218 73826 75454
rect 38382 75134 73826 75218
rect 38382 74898 46970 75134
rect 47206 74898 73826 75134
rect 74382 75218 77690 75454
rect 77926 75218 108410 75454
rect 108646 75218 109826 75454
rect 74382 75134 109826 75218
rect 74382 74898 77690 75134
rect 77926 74898 108410 75134
rect 108646 74898 109826 75134
rect 110382 75218 139130 75454
rect 139366 75218 145826 75454
rect 110382 75134 145826 75218
rect 110382 74898 139130 75134
rect 139366 74898 145826 75134
rect 146382 75218 169850 75454
rect 170086 75218 181826 75454
rect 146382 75134 181826 75218
rect 146382 74898 169850 75134
rect 170086 74898 181826 75134
rect 182382 75218 200570 75454
rect 200806 75218 217826 75454
rect 182382 75134 217826 75218
rect 182382 74898 200570 75134
rect 200806 74898 217826 75134
rect 218382 75218 231290 75454
rect 231526 75218 262010 75454
rect 262246 75218 289826 75454
rect 218382 75134 289826 75218
rect 218382 74898 231290 75134
rect 231526 74898 262010 75134
rect 262246 74898 289826 75134
rect 290382 74898 325826 75454
rect 326382 74898 361826 75454
rect 362382 74898 397826 75454
rect 398382 74898 433826 75454
rect 434382 74898 469826 75454
rect 470382 74898 505826 75454
rect 506382 74898 541826 75454
rect 542382 74898 577826 75454
rect 578382 74898 585342 75454
rect 585898 74898 592650 75454
rect -8726 74866 592650 74898
rect -8726 65494 592650 65526
rect -8726 64938 -8694 65494
rect -8138 64938 27866 65494
rect 28422 64938 63866 65494
rect 64422 64938 99866 65494
rect 100422 64938 135866 65494
rect 136422 64938 171866 65494
rect 172422 64938 243866 65494
rect 244422 64938 279866 65494
rect 280422 64938 315866 65494
rect 316422 64938 351866 65494
rect 352422 64938 387866 65494
rect 388422 64938 423866 65494
rect 424422 64938 459866 65494
rect 460422 64938 495866 65494
rect 496422 64938 531866 65494
rect 532422 64938 567866 65494
rect 568422 64938 592062 65494
rect 592618 64938 592650 65494
rect -8726 64906 592650 64938
rect -8726 61774 592650 61806
rect -8726 61218 -7734 61774
rect -7178 61218 60146 61774
rect 60702 61218 96146 61774
rect 96702 61218 132146 61774
rect 132702 61218 168146 61774
rect 168702 61218 204146 61774
rect 204702 61218 240146 61774
rect 240702 61218 276146 61774
rect 276702 61218 312146 61774
rect 312702 61218 348146 61774
rect 348702 61218 384146 61774
rect 384702 61218 420146 61774
rect 420702 61218 456146 61774
rect 456702 61218 492146 61774
rect 492702 61218 528146 61774
rect 528702 61218 564146 61774
rect 564702 61218 591102 61774
rect 591658 61218 592650 61774
rect -8726 61186 592650 61218
rect -8726 58054 592650 58086
rect -8726 57498 -6774 58054
rect -6218 57498 20426 58054
rect 20982 57818 39290 58054
rect 39526 57818 56426 58054
rect 20982 57734 56426 57818
rect 20982 57498 39290 57734
rect 39526 57498 56426 57734
rect 56982 57818 70010 58054
rect 70246 57818 100730 58054
rect 100966 57818 128426 58054
rect 56982 57734 128426 57818
rect 56982 57498 70010 57734
rect 70246 57498 100730 57734
rect 100966 57498 128426 57734
rect 128982 57818 131450 58054
rect 131686 57818 162170 58054
rect 162406 57818 164426 58054
rect 128982 57734 164426 57818
rect 128982 57498 131450 57734
rect 131686 57498 162170 57734
rect 162406 57498 164426 57734
rect 164982 57818 192890 58054
rect 193126 57818 223610 58054
rect 223846 57818 236426 58054
rect 164982 57734 236426 57818
rect 164982 57498 192890 57734
rect 193126 57498 223610 57734
rect 223846 57498 236426 57734
rect 236982 57818 254330 58054
rect 254566 57818 272426 58054
rect 236982 57734 272426 57818
rect 236982 57498 254330 57734
rect 254566 57498 272426 57734
rect 272982 57818 285050 58054
rect 285286 57818 308426 58054
rect 272982 57734 308426 57818
rect 272982 57498 285050 57734
rect 285286 57498 308426 57734
rect 308982 57498 344426 58054
rect 344982 57498 380426 58054
rect 380982 57498 416426 58054
rect 416982 57498 452426 58054
rect 452982 57498 488426 58054
rect 488982 57498 524426 58054
rect 524982 57498 560426 58054
rect 560982 57498 590142 58054
rect 590698 57498 592650 58054
rect -8726 57466 592650 57498
rect -8726 54334 592650 54366
rect -8726 53778 -5814 54334
rect -5258 54098 31610 54334
rect 31846 54098 52706 54334
rect -5258 54014 52706 54098
rect -5258 53778 31610 54014
rect 31846 53778 52706 54014
rect 53262 54098 62330 54334
rect 62566 54098 88706 54334
rect 53262 54014 88706 54098
rect 53262 53778 62330 54014
rect 62566 53778 88706 54014
rect 89262 54098 93050 54334
rect 93286 54098 123770 54334
rect 124006 54098 124706 54334
rect 89262 54014 124706 54098
rect 89262 53778 93050 54014
rect 93286 53778 123770 54014
rect 124006 53778 124706 54014
rect 125262 54098 154490 54334
rect 154726 54098 160706 54334
rect 125262 54014 160706 54098
rect 125262 53778 154490 54014
rect 154726 53778 160706 54014
rect 161262 54098 185210 54334
rect 185446 54098 196706 54334
rect 161262 54014 196706 54098
rect 161262 53778 185210 54014
rect 185446 53778 196706 54014
rect 197262 54098 215930 54334
rect 216166 54098 232706 54334
rect 197262 54014 232706 54098
rect 197262 53778 215930 54014
rect 216166 53778 232706 54014
rect 233262 54098 246650 54334
rect 246886 54098 268706 54334
rect 233262 54014 268706 54098
rect 233262 53778 246650 54014
rect 246886 53778 268706 54014
rect 269262 54098 277370 54334
rect 277606 54098 304706 54334
rect 269262 54014 304706 54098
rect 269262 53778 277370 54014
rect 277606 53778 304706 54014
rect 305262 53778 340706 54334
rect 341262 53778 376706 54334
rect 377262 53778 412706 54334
rect 413262 53778 448706 54334
rect 449262 53778 484706 54334
rect 485262 53778 520706 54334
rect 521262 53778 556706 54334
rect 557262 53778 589182 54334
rect 589738 53778 592650 54334
rect -8726 53746 592650 53778
rect -8726 50614 592650 50646
rect -8726 50058 -4854 50614
rect -4298 50058 12986 50614
rect 13542 50058 48986 50614
rect 49542 50058 120986 50614
rect 121542 50058 156986 50614
rect 157542 50058 228986 50614
rect 229542 50058 264986 50614
rect 265542 50058 300986 50614
rect 301542 50058 336986 50614
rect 337542 50058 372986 50614
rect 373542 50058 408986 50614
rect 409542 50058 444986 50614
rect 445542 50058 480986 50614
rect 481542 50058 516986 50614
rect 517542 50058 552986 50614
rect 553542 50058 588222 50614
rect 588778 50058 592650 50614
rect -8726 50026 592650 50058
rect -8726 46894 592650 46926
rect -8726 46338 -3894 46894
rect -3338 46338 9266 46894
rect 9822 46338 45266 46894
rect 45822 46338 81266 46894
rect 81822 46338 117266 46894
rect 117822 46338 153266 46894
rect 153822 46338 189266 46894
rect 189822 46338 225266 46894
rect 225822 46338 297266 46894
rect 297822 46338 333266 46894
rect 333822 46338 369266 46894
rect 369822 46338 405266 46894
rect 405822 46338 441266 46894
rect 441822 46338 477266 46894
rect 477822 46338 513266 46894
rect 513822 46338 549266 46894
rect 549822 46338 587262 46894
rect 587818 46338 592650 46894
rect -8726 46306 592650 46338
rect -8726 43174 592650 43206
rect -8726 42618 -2934 43174
rect -2378 42618 5546 43174
rect 6102 42938 17310 43174
rect 17546 42938 23930 43174
rect 24166 42938 41546 43174
rect 6102 42854 41546 42938
rect 6102 42618 17310 42854
rect 17546 42618 23930 42854
rect 24166 42618 41546 42854
rect 42102 42938 54650 43174
rect 54886 42938 85370 43174
rect 85606 42938 116090 43174
rect 116326 42938 146810 43174
rect 147046 42938 149546 43174
rect 42102 42854 149546 42938
rect 42102 42618 54650 42854
rect 54886 42618 85370 42854
rect 85606 42618 116090 42854
rect 116326 42618 146810 42854
rect 147046 42618 149546 42854
rect 150102 42938 177530 43174
rect 177766 42938 208250 43174
rect 208486 42938 221546 43174
rect 150102 42854 221546 42938
rect 150102 42618 177530 42854
rect 177766 42618 208250 42854
rect 208486 42618 221546 42854
rect 222102 42938 238970 43174
rect 239206 42938 257546 43174
rect 222102 42854 257546 42938
rect 222102 42618 238970 42854
rect 239206 42618 257546 42854
rect 258102 42938 269690 43174
rect 269926 42938 293546 43174
rect 258102 42854 293546 42938
rect 258102 42618 269690 42854
rect 269926 42618 293546 42854
rect 294102 42618 329546 43174
rect 330102 42618 365546 43174
rect 366102 42618 401546 43174
rect 402102 42618 437546 43174
rect 438102 42618 473546 43174
rect 474102 42618 509546 43174
rect 510102 42618 545546 43174
rect 546102 42618 581546 43174
rect 582102 42618 586302 43174
rect 586858 42618 592650 43174
rect -8726 42586 592650 42618
rect -8726 39454 592650 39486
rect -8726 38898 -1974 39454
rect -1418 38898 1826 39454
rect 2382 39218 16250 39454
rect 16486 39218 37826 39454
rect 2382 39134 37826 39218
rect 2382 38898 16250 39134
rect 16486 38898 37826 39134
rect 38382 39218 46970 39454
rect 47206 39218 73826 39454
rect 38382 39134 73826 39218
rect 38382 38898 46970 39134
rect 47206 38898 73826 39134
rect 74382 39218 77690 39454
rect 77926 39218 108410 39454
rect 108646 39218 109826 39454
rect 74382 39134 109826 39218
rect 74382 38898 77690 39134
rect 77926 38898 108410 39134
rect 108646 38898 109826 39134
rect 110382 39218 139130 39454
rect 139366 39218 145826 39454
rect 110382 39134 145826 39218
rect 110382 38898 139130 39134
rect 139366 38898 145826 39134
rect 146382 39218 169850 39454
rect 170086 39218 181826 39454
rect 146382 39134 181826 39218
rect 146382 38898 169850 39134
rect 170086 38898 181826 39134
rect 182382 39218 200570 39454
rect 200806 39218 217826 39454
rect 182382 39134 217826 39218
rect 182382 38898 200570 39134
rect 200806 38898 217826 39134
rect 218382 39218 231290 39454
rect 231526 39218 262010 39454
rect 262246 39218 289826 39454
rect 218382 39134 289826 39218
rect 218382 38898 231290 39134
rect 231526 38898 262010 39134
rect 262246 38898 289826 39134
rect 290382 38898 325826 39454
rect 326382 38898 361826 39454
rect 362382 38898 397826 39454
rect 398382 38898 433826 39454
rect 434382 38898 469826 39454
rect 470382 38898 505826 39454
rect 506382 38898 541826 39454
rect 542382 38898 577826 39454
rect 578382 38898 585342 39454
rect 585898 38898 592650 39454
rect -8726 38866 592650 38898
rect -8726 29494 592650 29526
rect -8726 28938 -8694 29494
rect -8138 28938 27866 29494
rect 28422 28938 63866 29494
rect 64422 28938 99866 29494
rect 100422 28938 135866 29494
rect 136422 28938 171866 29494
rect 172422 28938 243866 29494
rect 244422 28938 279866 29494
rect 280422 28938 315866 29494
rect 316422 28938 351866 29494
rect 352422 28938 387866 29494
rect 388422 28938 423866 29494
rect 424422 28938 459866 29494
rect 460422 28938 495866 29494
rect 496422 28938 531866 29494
rect 532422 28938 567866 29494
rect 568422 28938 592062 29494
rect 592618 28938 592650 29494
rect -8726 28906 592650 28938
rect -8726 25774 592650 25806
rect -8726 25218 -7734 25774
rect -7178 25218 60146 25774
rect 60702 25218 96146 25774
rect 96702 25218 132146 25774
rect 132702 25218 168146 25774
rect 168702 25218 204146 25774
rect 204702 25218 240146 25774
rect 240702 25218 276146 25774
rect 276702 25218 312146 25774
rect 312702 25218 348146 25774
rect 348702 25218 384146 25774
rect 384702 25218 420146 25774
rect 420702 25218 456146 25774
rect 456702 25218 492146 25774
rect 492702 25218 528146 25774
rect 528702 25218 564146 25774
rect 564702 25218 591102 25774
rect 591658 25218 592650 25774
rect -8726 25186 592650 25218
rect -8726 22054 592650 22086
rect -8726 21498 -6774 22054
rect -6218 21498 20426 22054
rect 20982 21818 39290 22054
rect 39526 21818 56426 22054
rect 20982 21734 56426 21818
rect 20982 21498 39290 21734
rect 39526 21498 56426 21734
rect 56982 21818 70010 22054
rect 70246 21818 100730 22054
rect 100966 21818 128426 22054
rect 56982 21734 128426 21818
rect 56982 21498 70010 21734
rect 70246 21498 100730 21734
rect 100966 21498 128426 21734
rect 128982 21818 131450 22054
rect 131686 21818 162170 22054
rect 162406 21818 164426 22054
rect 128982 21734 164426 21818
rect 128982 21498 131450 21734
rect 131686 21498 162170 21734
rect 162406 21498 164426 21734
rect 164982 21818 192890 22054
rect 193126 21818 223610 22054
rect 223846 21818 236426 22054
rect 164982 21734 236426 21818
rect 164982 21498 192890 21734
rect 193126 21498 223610 21734
rect 223846 21498 236426 21734
rect 236982 21818 254330 22054
rect 254566 21818 272426 22054
rect 236982 21734 272426 21818
rect 236982 21498 254330 21734
rect 254566 21498 272426 21734
rect 272982 21818 285050 22054
rect 285286 21818 308426 22054
rect 272982 21734 308426 21818
rect 272982 21498 285050 21734
rect 285286 21498 308426 21734
rect 308982 21498 344426 22054
rect 344982 21498 380426 22054
rect 380982 21498 416426 22054
rect 416982 21498 452426 22054
rect 452982 21498 488426 22054
rect 488982 21498 524426 22054
rect 524982 21498 560426 22054
rect 560982 21498 590142 22054
rect 590698 21498 592650 22054
rect -8726 21466 592650 21498
rect -8726 18334 592650 18366
rect -8726 17778 -5814 18334
rect -5258 18098 31610 18334
rect 31846 18098 52706 18334
rect -5258 18014 52706 18098
rect -5258 17778 31610 18014
rect 31846 17778 52706 18014
rect 53262 18098 62330 18334
rect 62566 18098 88706 18334
rect 53262 18014 88706 18098
rect 53262 17778 62330 18014
rect 62566 17778 88706 18014
rect 89262 18098 93050 18334
rect 93286 18098 123770 18334
rect 124006 18098 124706 18334
rect 89262 18014 124706 18098
rect 89262 17778 93050 18014
rect 93286 17778 123770 18014
rect 124006 17778 124706 18014
rect 125262 18098 154490 18334
rect 154726 18098 160706 18334
rect 125262 18014 160706 18098
rect 125262 17778 154490 18014
rect 154726 17778 160706 18014
rect 161262 18098 185210 18334
rect 185446 18098 196706 18334
rect 161262 18014 196706 18098
rect 161262 17778 185210 18014
rect 185446 17778 196706 18014
rect 197262 18098 215930 18334
rect 216166 18098 232706 18334
rect 197262 18014 232706 18098
rect 197262 17778 215930 18014
rect 216166 17778 232706 18014
rect 233262 18098 246650 18334
rect 246886 18098 268706 18334
rect 233262 18014 268706 18098
rect 233262 17778 246650 18014
rect 246886 17778 268706 18014
rect 269262 18098 277370 18334
rect 277606 18098 304706 18334
rect 269262 18014 304706 18098
rect 269262 17778 277370 18014
rect 277606 17778 304706 18014
rect 305262 17778 340706 18334
rect 341262 17778 376706 18334
rect 377262 17778 412706 18334
rect 413262 17778 448706 18334
rect 449262 17778 484706 18334
rect 485262 17778 520706 18334
rect 521262 17778 556706 18334
rect 557262 17778 589182 18334
rect 589738 17778 592650 18334
rect -8726 17746 592650 17778
rect -8726 14614 592650 14646
rect -8726 14058 -4854 14614
rect -4298 14058 12986 14614
rect 13542 14058 48986 14614
rect 49542 14058 120986 14614
rect 121542 14058 156986 14614
rect 157542 14058 228986 14614
rect 229542 14058 264986 14614
rect 265542 14058 300986 14614
rect 301542 14058 336986 14614
rect 337542 14058 372986 14614
rect 373542 14058 408986 14614
rect 409542 14058 444986 14614
rect 445542 14058 480986 14614
rect 481542 14058 516986 14614
rect 517542 14058 552986 14614
rect 553542 14058 588222 14614
rect 588778 14058 592650 14614
rect -8726 14026 592650 14058
rect -8726 10894 592650 10926
rect -8726 10338 -3894 10894
rect -3338 10338 9266 10894
rect 9822 10338 45266 10894
rect 45822 10338 81266 10894
rect 81822 10338 117266 10894
rect 117822 10338 153266 10894
rect 153822 10338 189266 10894
rect 189822 10338 225266 10894
rect 225822 10338 297266 10894
rect 297822 10338 333266 10894
rect 333822 10338 369266 10894
rect 369822 10338 405266 10894
rect 405822 10338 441266 10894
rect 441822 10338 477266 10894
rect 477822 10338 513266 10894
rect 513822 10338 549266 10894
rect 549822 10338 587262 10894
rect 587818 10338 592650 10894
rect -8726 10306 592650 10338
rect -8726 7174 592650 7206
rect -8726 6618 -2934 7174
rect -2378 6618 5546 7174
rect 6102 6938 17310 7174
rect 17546 6938 23930 7174
rect 24166 6938 41546 7174
rect 6102 6854 41546 6938
rect 6102 6618 17310 6854
rect 17546 6618 23930 6854
rect 24166 6618 41546 6854
rect 42102 6938 54650 7174
rect 54886 6938 85370 7174
rect 85606 6938 116090 7174
rect 116326 6938 146810 7174
rect 147046 6938 149546 7174
rect 42102 6854 149546 6938
rect 42102 6618 54650 6854
rect 54886 6618 85370 6854
rect 85606 6618 116090 6854
rect 116326 6618 146810 6854
rect 147046 6618 149546 6854
rect 150102 6938 177530 7174
rect 177766 6938 208250 7174
rect 208486 6938 221546 7174
rect 150102 6854 221546 6938
rect 150102 6618 177530 6854
rect 177766 6618 208250 6854
rect 208486 6618 221546 6854
rect 222102 6938 238970 7174
rect 239206 6938 257546 7174
rect 222102 6854 257546 6938
rect 222102 6618 238970 6854
rect 239206 6618 257546 6854
rect 258102 6938 269690 7174
rect 269926 6938 293546 7174
rect 258102 6854 293546 6938
rect 258102 6618 269690 6854
rect 269926 6618 293546 6854
rect 294102 6618 329546 7174
rect 330102 6618 365546 7174
rect 366102 6618 401546 7174
rect 402102 6618 437546 7174
rect 438102 6618 473546 7174
rect 474102 6618 509546 7174
rect 510102 6618 545546 7174
rect 546102 6618 581546 7174
rect 582102 6618 586302 7174
rect 586858 6618 592650 7174
rect -8726 6586 592650 6618
rect -8726 3454 592650 3486
rect -8726 2898 -1974 3454
rect -1418 2898 1826 3454
rect 2382 2898 37826 3454
rect 38382 2898 73826 3454
rect 74382 2898 109826 3454
rect 110382 2898 145826 3454
rect 146382 2898 181826 3454
rect 182382 2898 217826 3454
rect 218382 2898 289826 3454
rect 290382 2898 325826 3454
rect 326382 2898 361826 3454
rect 362382 2898 397826 3454
rect 398382 2898 433826 3454
rect 434382 2898 469826 3454
rect 470382 2898 505826 3454
rect 506382 2898 541826 3454
rect 542382 2898 577826 3454
rect 578382 2898 585342 3454
rect 585898 2898 592650 3454
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -902 -1974 -346
rect -1418 -902 1826 -346
rect 2382 -902 37826 -346
rect 38382 -902 73826 -346
rect 74382 -902 109826 -346
rect 110382 -902 145826 -346
rect 146382 -902 181826 -346
rect 182382 -902 217826 -346
rect 218382 -902 253826 -346
rect 254382 -902 289826 -346
rect 290382 -902 325826 -346
rect 326382 -902 361826 -346
rect 362382 -902 397826 -346
rect 398382 -902 433826 -346
rect 434382 -902 469826 -346
rect 470382 -902 505826 -346
rect 506382 -902 541826 -346
rect 542382 -902 577826 -346
rect 578382 -902 585342 -346
rect 585898 -902 585930 -346
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1862 -2934 -1306
rect -2378 -1862 5546 -1306
rect 6102 -1862 41546 -1306
rect 42102 -1862 77546 -1306
rect 78102 -1862 113546 -1306
rect 114102 -1862 149546 -1306
rect 150102 -1862 185546 -1306
rect 186102 -1862 221546 -1306
rect 222102 -1862 257546 -1306
rect 258102 -1862 293546 -1306
rect 294102 -1862 329546 -1306
rect 330102 -1862 365546 -1306
rect 366102 -1862 401546 -1306
rect 402102 -1862 437546 -1306
rect 438102 -1862 473546 -1306
rect 474102 -1862 509546 -1306
rect 510102 -1862 545546 -1306
rect 546102 -1862 581546 -1306
rect 582102 -1862 586302 -1306
rect 586858 -1862 586890 -1306
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2822 -3894 -2266
rect -3338 -2822 9266 -2266
rect 9822 -2822 45266 -2266
rect 45822 -2822 81266 -2266
rect 81822 -2822 117266 -2266
rect 117822 -2822 153266 -2266
rect 153822 -2822 189266 -2266
rect 189822 -2822 225266 -2266
rect 225822 -2822 261266 -2266
rect 261822 -2822 297266 -2266
rect 297822 -2822 333266 -2266
rect 333822 -2822 369266 -2266
rect 369822 -2822 405266 -2266
rect 405822 -2822 441266 -2266
rect 441822 -2822 477266 -2266
rect 477822 -2822 513266 -2266
rect 513822 -2822 549266 -2266
rect 549822 -2822 587262 -2266
rect 587818 -2822 587850 -2266
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3782 -4854 -3226
rect -4298 -3782 12986 -3226
rect 13542 -3782 48986 -3226
rect 49542 -3782 84986 -3226
rect 85542 -3782 120986 -3226
rect 121542 -3782 156986 -3226
rect 157542 -3782 192986 -3226
rect 193542 -3782 228986 -3226
rect 229542 -3782 264986 -3226
rect 265542 -3782 300986 -3226
rect 301542 -3782 336986 -3226
rect 337542 -3782 372986 -3226
rect 373542 -3782 408986 -3226
rect 409542 -3782 444986 -3226
rect 445542 -3782 480986 -3226
rect 481542 -3782 516986 -3226
rect 517542 -3782 552986 -3226
rect 553542 -3782 588222 -3226
rect 588778 -3782 588810 -3226
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4742 -5814 -4186
rect -5258 -4742 16706 -4186
rect 17262 -4742 52706 -4186
rect 53262 -4742 88706 -4186
rect 89262 -4742 124706 -4186
rect 125262 -4742 160706 -4186
rect 161262 -4742 196706 -4186
rect 197262 -4742 232706 -4186
rect 233262 -4742 268706 -4186
rect 269262 -4742 304706 -4186
rect 305262 -4742 340706 -4186
rect 341262 -4742 376706 -4186
rect 377262 -4742 412706 -4186
rect 413262 -4742 448706 -4186
rect 449262 -4742 484706 -4186
rect 485262 -4742 520706 -4186
rect 521262 -4742 556706 -4186
rect 557262 -4742 589182 -4186
rect 589738 -4742 589770 -4186
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5702 -6774 -5146
rect -6218 -5702 20426 -5146
rect 20982 -5702 56426 -5146
rect 56982 -5702 92426 -5146
rect 92982 -5702 128426 -5146
rect 128982 -5702 164426 -5146
rect 164982 -5702 200426 -5146
rect 200982 -5702 236426 -5146
rect 236982 -5702 272426 -5146
rect 272982 -5702 308426 -5146
rect 308982 -5702 344426 -5146
rect 344982 -5702 380426 -5146
rect 380982 -5702 416426 -5146
rect 416982 -5702 452426 -5146
rect 452982 -5702 488426 -5146
rect 488982 -5702 524426 -5146
rect 524982 -5702 560426 -5146
rect 560982 -5702 590142 -5146
rect 590698 -5702 590730 -5146
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6662 -7734 -6106
rect -7178 -6662 24146 -6106
rect 24702 -6662 60146 -6106
rect 60702 -6662 96146 -6106
rect 96702 -6662 132146 -6106
rect 132702 -6662 168146 -6106
rect 168702 -6662 204146 -6106
rect 204702 -6662 240146 -6106
rect 240702 -6662 276146 -6106
rect 276702 -6662 312146 -6106
rect 312702 -6662 348146 -6106
rect 348702 -6662 384146 -6106
rect 384702 -6662 420146 -6106
rect 420702 -6662 456146 -6106
rect 456702 -6662 492146 -6106
rect 492702 -6662 528146 -6106
rect 528702 -6662 564146 -6106
rect 564702 -6662 591102 -6106
rect 591658 -6662 591690 -6106
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7622 -8694 -7066
rect -8138 -7622 27866 -7066
rect 28422 -7622 63866 -7066
rect 64422 -7622 99866 -7066
rect 100422 -7622 135866 -7066
rect 136422 -7622 171866 -7066
rect 172422 -7622 207866 -7066
rect 208422 -7622 243866 -7066
rect 244422 -7622 279866 -7066
rect 280422 -7622 315866 -7066
rect 316422 -7622 351866 -7066
rect 352422 -7622 387866 -7066
rect 388422 -7622 423866 -7066
rect 424422 -7622 459866 -7066
rect 460422 -7622 495866 -7066
rect 496422 -7622 531866 -7066
rect 532422 -7622 567866 -7066
rect 568422 -7622 592062 -7066
rect 592618 -7622 592650 -7066
rect -8726 -7654 592650 -7622
use user_proj_example  mprj
timestamp 0
transform 1 0 12000 0 1 3000
box 0 0 278890 277488
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 1200 0 0 0 analog_io[0]
port 1 nsew
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 560 90 0 0 analog_io[10]
port 2 nsew
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 560 90 0 0 analog_io[11]
port 3 nsew
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 560 90 0 0 analog_io[12]
port 4 nsew
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 560 90 0 0 analog_io[13]
port 5 nsew
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 560 90 0 0 analog_io[14]
port 6 nsew
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 560 90 0 0 analog_io[15]
port 7 nsew
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 560 90 0 0 analog_io[16]
port 8 nsew
flabel metal3 s -960 697220 480 697460 0 FreeSans 1200 0 0 0 analog_io[17]
port 9 nsew
flabel metal3 s -960 644996 480 645236 0 FreeSans 1200 0 0 0 analog_io[18]
port 10 nsew
flabel metal3 s -960 592908 480 593148 0 FreeSans 1200 0 0 0 analog_io[19]
port 11 nsew
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 1200 0 0 0 analog_io[1]
port 12 nsew
flabel metal3 s -960 540684 480 540924 0 FreeSans 1200 0 0 0 analog_io[20]
port 13 nsew
flabel metal3 s -960 488596 480 488836 0 FreeSans 1200 0 0 0 analog_io[21]
port 14 nsew
flabel metal3 s -960 436508 480 436748 0 FreeSans 1200 0 0 0 analog_io[22]
port 15 nsew
flabel metal3 s -960 384284 480 384524 0 FreeSans 1200 0 0 0 analog_io[23]
port 16 nsew
flabel metal3 s -960 332196 480 332436 0 FreeSans 1200 0 0 0 analog_io[24]
port 17 nsew
flabel metal3 s -960 279972 480 280212 0 FreeSans 1200 0 0 0 analog_io[25]
port 18 nsew
flabel metal3 s -960 227884 480 228124 0 FreeSans 1200 0 0 0 analog_io[26]
port 19 nsew
flabel metal3 s -960 175796 480 176036 0 FreeSans 1200 0 0 0 analog_io[27]
port 20 nsew
flabel metal3 s -960 123572 480 123812 0 FreeSans 1200 0 0 0 analog_io[28]
port 21 nsew
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 1200 0 0 0 analog_io[2]
port 22 nsew
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 1200 0 0 0 analog_io[3]
port 23 nsew
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 1200 0 0 0 analog_io[4]
port 24 nsew
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 1200 0 0 0 analog_io[5]
port 25 nsew
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 1200 0 0 0 analog_io[6]
port 26 nsew
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 1200 0 0 0 analog_io[7]
port 27 nsew
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 560 90 0 0 analog_io[8]
port 28 nsew
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 560 90 0 0 analog_io[9]
port 29 nsew
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 1200 0 0 0 io_in[0]
port 30 nsew
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 1200 0 0 0 io_in[10]
port 31 nsew
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 1200 0 0 0 io_in[11]
port 32 nsew
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 1200 0 0 0 io_in[12]
port 33 nsew
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 1200 0 0 0 io_in[13]
port 34 nsew
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 1200 0 0 0 io_in[14]
port 35 nsew
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 560 90 0 0 io_in[15]
port 36 nsew
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 560 90 0 0 io_in[16]
port 37 nsew
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 560 90 0 0 io_in[17]
port 38 nsew
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 560 90 0 0 io_in[18]
port 39 nsew
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 560 90 0 0 io_in[19]
port 40 nsew
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 1200 0 0 0 io_in[1]
port 41 nsew
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 560 90 0 0 io_in[20]
port 42 nsew
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 560 90 0 0 io_in[21]
port 43 nsew
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 560 90 0 0 io_in[22]
port 44 nsew
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 560 90 0 0 io_in[23]
port 45 nsew
flabel metal3 s -960 684164 480 684404 0 FreeSans 1200 0 0 0 io_in[24]
port 46 nsew
flabel metal3 s -960 631940 480 632180 0 FreeSans 1200 0 0 0 io_in[25]
port 47 nsew
flabel metal3 s -960 579852 480 580092 0 FreeSans 1200 0 0 0 io_in[26]
port 48 nsew
flabel metal3 s -960 527764 480 528004 0 FreeSans 1200 0 0 0 io_in[27]
port 49 nsew
flabel metal3 s -960 475540 480 475780 0 FreeSans 1200 0 0 0 io_in[28]
port 50 nsew
flabel metal3 s -960 423452 480 423692 0 FreeSans 1200 0 0 0 io_in[29]
port 51 nsew
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 1200 0 0 0 io_in[2]
port 52 nsew
flabel metal3 s -960 371228 480 371468 0 FreeSans 1200 0 0 0 io_in[30]
port 53 nsew
flabel metal3 s -960 319140 480 319380 0 FreeSans 1200 0 0 0 io_in[31]
port 54 nsew
flabel metal3 s -960 267052 480 267292 0 FreeSans 1200 0 0 0 io_in[32]
port 55 nsew
flabel metal3 s -960 214828 480 215068 0 FreeSans 1200 0 0 0 io_in[33]
port 56 nsew
flabel metal3 s -960 162740 480 162980 0 FreeSans 1200 0 0 0 io_in[34]
port 57 nsew
flabel metal3 s -960 110516 480 110756 0 FreeSans 1200 0 0 0 io_in[35]
port 58 nsew
flabel metal3 s -960 71484 480 71724 0 FreeSans 1200 0 0 0 io_in[36]
port 59 nsew
flabel metal3 s -960 32316 480 32556 0 FreeSans 1200 0 0 0 io_in[37]
port 60 nsew
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 1200 0 0 0 io_in[3]
port 61 nsew
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 1200 0 0 0 io_in[4]
port 62 nsew
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 1200 0 0 0 io_in[5]
port 63 nsew
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 1200 0 0 0 io_in[6]
port 64 nsew
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 1200 0 0 0 io_in[7]
port 65 nsew
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 1200 0 0 0 io_in[8]
port 66 nsew
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 1200 0 0 0 io_in[9]
port 67 nsew
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 1200 0 0 0 io_oeb[0]
port 68 nsew
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 1200 0 0 0 io_oeb[10]
port 69 nsew
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 1200 0 0 0 io_oeb[11]
port 70 nsew
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 1200 0 0 0 io_oeb[12]
port 71 nsew
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 1200 0 0 0 io_oeb[13]
port 72 nsew
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 1200 0 0 0 io_oeb[14]
port 73 nsew
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 560 90 0 0 io_oeb[15]
port 74 nsew
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 560 90 0 0 io_oeb[16]
port 75 nsew
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 560 90 0 0 io_oeb[17]
port 76 nsew
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 560 90 0 0 io_oeb[18]
port 77 nsew
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 560 90 0 0 io_oeb[19]
port 78 nsew
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 1200 0 0 0 io_oeb[1]
port 79 nsew
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 560 90 0 0 io_oeb[20]
port 80 nsew
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 560 90 0 0 io_oeb[21]
port 81 nsew
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 560 90 0 0 io_oeb[22]
port 82 nsew
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 560 90 0 0 io_oeb[23]
port 83 nsew
flabel metal3 s -960 658052 480 658292 0 FreeSans 1200 0 0 0 io_oeb[24]
port 84 nsew
flabel metal3 s -960 605964 480 606204 0 FreeSans 1200 0 0 0 io_oeb[25]
port 85 nsew
flabel metal3 s -960 553740 480 553980 0 FreeSans 1200 0 0 0 io_oeb[26]
port 86 nsew
flabel metal3 s -960 501652 480 501892 0 FreeSans 1200 0 0 0 io_oeb[27]
port 87 nsew
flabel metal3 s -960 449428 480 449668 0 FreeSans 1200 0 0 0 io_oeb[28]
port 88 nsew
flabel metal3 s -960 397340 480 397580 0 FreeSans 1200 0 0 0 io_oeb[29]
port 89 nsew
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 1200 0 0 0 io_oeb[2]
port 90 nsew
flabel metal3 s -960 345252 480 345492 0 FreeSans 1200 0 0 0 io_oeb[30]
port 91 nsew
flabel metal3 s -960 293028 480 293268 0 FreeSans 1200 0 0 0 io_oeb[31]
port 92 nsew
flabel metal3 s -960 240940 480 241180 0 FreeSans 1200 0 0 0 io_oeb[32]
port 93 nsew
flabel metal3 s -960 188716 480 188956 0 FreeSans 1200 0 0 0 io_oeb[33]
port 94 nsew
flabel metal3 s -960 136628 480 136868 0 FreeSans 1200 0 0 0 io_oeb[34]
port 95 nsew
flabel metal3 s -960 84540 480 84780 0 FreeSans 1200 0 0 0 io_oeb[35]
port 96 nsew
flabel metal3 s -960 45372 480 45612 0 FreeSans 1200 0 0 0 io_oeb[36]
port 97 nsew
flabel metal3 s -960 6340 480 6580 0 FreeSans 1200 0 0 0 io_oeb[37]
port 98 nsew
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 1200 0 0 0 io_oeb[3]
port 99 nsew
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 1200 0 0 0 io_oeb[4]
port 100 nsew
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 1200 0 0 0 io_oeb[5]
port 101 nsew
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 1200 0 0 0 io_oeb[6]
port 102 nsew
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 1200 0 0 0 io_oeb[7]
port 103 nsew
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 1200 0 0 0 io_oeb[8]
port 104 nsew
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 1200 0 0 0 io_oeb[9]
port 105 nsew
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 1200 0 0 0 io_out[0]
port 106 nsew
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 1200 0 0 0 io_out[10]
port 107 nsew
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 1200 0 0 0 io_out[11]
port 108 nsew
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 1200 0 0 0 io_out[12]
port 109 nsew
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 1200 0 0 0 io_out[13]
port 110 nsew
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 1200 0 0 0 io_out[14]
port 111 nsew
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 560 90 0 0 io_out[15]
port 112 nsew
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 560 90 0 0 io_out[16]
port 113 nsew
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 560 90 0 0 io_out[17]
port 114 nsew
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 560 90 0 0 io_out[18]
port 115 nsew
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 560 90 0 0 io_out[19]
port 116 nsew
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 1200 0 0 0 io_out[1]
port 117 nsew
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 560 90 0 0 io_out[20]
port 118 nsew
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 560 90 0 0 io_out[21]
port 119 nsew
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 560 90 0 0 io_out[22]
port 120 nsew
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 560 90 0 0 io_out[23]
port 121 nsew
flabel metal3 s -960 671108 480 671348 0 FreeSans 1200 0 0 0 io_out[24]
port 122 nsew
flabel metal3 s -960 619020 480 619260 0 FreeSans 1200 0 0 0 io_out[25]
port 123 nsew
flabel metal3 s -960 566796 480 567036 0 FreeSans 1200 0 0 0 io_out[26]
port 124 nsew
flabel metal3 s -960 514708 480 514948 0 FreeSans 1200 0 0 0 io_out[27]
port 125 nsew
flabel metal3 s -960 462484 480 462724 0 FreeSans 1200 0 0 0 io_out[28]
port 126 nsew
flabel metal3 s -960 410396 480 410636 0 FreeSans 1200 0 0 0 io_out[29]
port 127 nsew
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 1200 0 0 0 io_out[2]
port 128 nsew
flabel metal3 s -960 358308 480 358548 0 FreeSans 1200 0 0 0 io_out[30]
port 129 nsew
flabel metal3 s -960 306084 480 306324 0 FreeSans 1200 0 0 0 io_out[31]
port 130 nsew
flabel metal3 s -960 253996 480 254236 0 FreeSans 1200 0 0 0 io_out[32]
port 131 nsew
flabel metal3 s -960 201772 480 202012 0 FreeSans 1200 0 0 0 io_out[33]
port 132 nsew
flabel metal3 s -960 149684 480 149924 0 FreeSans 1200 0 0 0 io_out[34]
port 133 nsew
flabel metal3 s -960 97460 480 97700 0 FreeSans 1200 0 0 0 io_out[35]
port 134 nsew
flabel metal3 s -960 58428 480 58668 0 FreeSans 1200 0 0 0 io_out[36]
port 135 nsew
flabel metal3 s -960 19260 480 19500 0 FreeSans 1200 0 0 0 io_out[37]
port 136 nsew
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 1200 0 0 0 io_out[3]
port 137 nsew
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 1200 0 0 0 io_out[4]
port 138 nsew
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 1200 0 0 0 io_out[5]
port 139 nsew
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 1200 0 0 0 io_out[6]
port 140 nsew
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 1200 0 0 0 io_out[7]
port 141 nsew
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 1200 0 0 0 io_out[8]
port 142 nsew
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 1200 0 0 0 io_out[9]
port 143 nsew
flabel metal2 s 125846 -960 125958 480 0 FreeSans 560 90 0 0 la_data_in[0]
port 144 nsew
flabel metal2 s 480506 -960 480618 480 0 FreeSans 560 90 0 0 la_data_in[100]
port 145 nsew
flabel metal2 s 484002 -960 484114 480 0 FreeSans 560 90 0 0 la_data_in[101]
port 146 nsew
flabel metal2 s 487590 -960 487702 480 0 FreeSans 560 90 0 0 la_data_in[102]
port 147 nsew
flabel metal2 s 491086 -960 491198 480 0 FreeSans 560 90 0 0 la_data_in[103]
port 148 nsew
flabel metal2 s 494674 -960 494786 480 0 FreeSans 560 90 0 0 la_data_in[104]
port 149 nsew
flabel metal2 s 498170 -960 498282 480 0 FreeSans 560 90 0 0 la_data_in[105]
port 150 nsew
flabel metal2 s 501758 -960 501870 480 0 FreeSans 560 90 0 0 la_data_in[106]
port 151 nsew
flabel metal2 s 505346 -960 505458 480 0 FreeSans 560 90 0 0 la_data_in[107]
port 152 nsew
flabel metal2 s 508842 -960 508954 480 0 FreeSans 560 90 0 0 la_data_in[108]
port 153 nsew
flabel metal2 s 512430 -960 512542 480 0 FreeSans 560 90 0 0 la_data_in[109]
port 154 nsew
flabel metal2 s 161266 -960 161378 480 0 FreeSans 560 90 0 0 la_data_in[10]
port 155 nsew
flabel metal2 s 515926 -960 516038 480 0 FreeSans 560 90 0 0 la_data_in[110]
port 156 nsew
flabel metal2 s 519514 -960 519626 480 0 FreeSans 560 90 0 0 la_data_in[111]
port 157 nsew
flabel metal2 s 523010 -960 523122 480 0 FreeSans 560 90 0 0 la_data_in[112]
port 158 nsew
flabel metal2 s 526598 -960 526710 480 0 FreeSans 560 90 0 0 la_data_in[113]
port 159 nsew
flabel metal2 s 530094 -960 530206 480 0 FreeSans 560 90 0 0 la_data_in[114]
port 160 nsew
flabel metal2 s 533682 -960 533794 480 0 FreeSans 560 90 0 0 la_data_in[115]
port 161 nsew
flabel metal2 s 537178 -960 537290 480 0 FreeSans 560 90 0 0 la_data_in[116]
port 162 nsew
flabel metal2 s 540766 -960 540878 480 0 FreeSans 560 90 0 0 la_data_in[117]
port 163 nsew
flabel metal2 s 544354 -960 544466 480 0 FreeSans 560 90 0 0 la_data_in[118]
port 164 nsew
flabel metal2 s 547850 -960 547962 480 0 FreeSans 560 90 0 0 la_data_in[119]
port 165 nsew
flabel metal2 s 164854 -960 164966 480 0 FreeSans 560 90 0 0 la_data_in[11]
port 166 nsew
flabel metal2 s 551438 -960 551550 480 0 FreeSans 560 90 0 0 la_data_in[120]
port 167 nsew
flabel metal2 s 554934 -960 555046 480 0 FreeSans 560 90 0 0 la_data_in[121]
port 168 nsew
flabel metal2 s 558522 -960 558634 480 0 FreeSans 560 90 0 0 la_data_in[122]
port 169 nsew
flabel metal2 s 562018 -960 562130 480 0 FreeSans 560 90 0 0 la_data_in[123]
port 170 nsew
flabel metal2 s 565606 -960 565718 480 0 FreeSans 560 90 0 0 la_data_in[124]
port 171 nsew
flabel metal2 s 569102 -960 569214 480 0 FreeSans 560 90 0 0 la_data_in[125]
port 172 nsew
flabel metal2 s 572690 -960 572802 480 0 FreeSans 560 90 0 0 la_data_in[126]
port 173 nsew
flabel metal2 s 576278 -960 576390 480 0 FreeSans 560 90 0 0 la_data_in[127]
port 174 nsew
flabel metal2 s 168350 -960 168462 480 0 FreeSans 560 90 0 0 la_data_in[12]
port 175 nsew
flabel metal2 s 171938 -960 172050 480 0 FreeSans 560 90 0 0 la_data_in[13]
port 176 nsew
flabel metal2 s 175434 -960 175546 480 0 FreeSans 560 90 0 0 la_data_in[14]
port 177 nsew
flabel metal2 s 179022 -960 179134 480 0 FreeSans 560 90 0 0 la_data_in[15]
port 178 nsew
flabel metal2 s 182518 -960 182630 480 0 FreeSans 560 90 0 0 la_data_in[16]
port 179 nsew
flabel metal2 s 186106 -960 186218 480 0 FreeSans 560 90 0 0 la_data_in[17]
port 180 nsew
flabel metal2 s 189694 -960 189806 480 0 FreeSans 560 90 0 0 la_data_in[18]
port 181 nsew
flabel metal2 s 193190 -960 193302 480 0 FreeSans 560 90 0 0 la_data_in[19]
port 182 nsew
flabel metal2 s 129342 -960 129454 480 0 FreeSans 560 90 0 0 la_data_in[1]
port 183 nsew
flabel metal2 s 196778 -960 196890 480 0 FreeSans 560 90 0 0 la_data_in[20]
port 184 nsew
flabel metal2 s 200274 -960 200386 480 0 FreeSans 560 90 0 0 la_data_in[21]
port 185 nsew
flabel metal2 s 203862 -960 203974 480 0 FreeSans 560 90 0 0 la_data_in[22]
port 186 nsew
flabel metal2 s 207358 -960 207470 480 0 FreeSans 560 90 0 0 la_data_in[23]
port 187 nsew
flabel metal2 s 210946 -960 211058 480 0 FreeSans 560 90 0 0 la_data_in[24]
port 188 nsew
flabel metal2 s 214442 -960 214554 480 0 FreeSans 560 90 0 0 la_data_in[25]
port 189 nsew
flabel metal2 s 218030 -960 218142 480 0 FreeSans 560 90 0 0 la_data_in[26]
port 190 nsew
flabel metal2 s 221526 -960 221638 480 0 FreeSans 560 90 0 0 la_data_in[27]
port 191 nsew
flabel metal2 s 225114 -960 225226 480 0 FreeSans 560 90 0 0 la_data_in[28]
port 192 nsew
flabel metal2 s 228702 -960 228814 480 0 FreeSans 560 90 0 0 la_data_in[29]
port 193 nsew
flabel metal2 s 132930 -960 133042 480 0 FreeSans 560 90 0 0 la_data_in[2]
port 194 nsew
flabel metal2 s 232198 -960 232310 480 0 FreeSans 560 90 0 0 la_data_in[30]
port 195 nsew
flabel metal2 s 235786 -960 235898 480 0 FreeSans 560 90 0 0 la_data_in[31]
port 196 nsew
flabel metal2 s 239282 -960 239394 480 0 FreeSans 560 90 0 0 la_data_in[32]
port 197 nsew
flabel metal2 s 242870 -960 242982 480 0 FreeSans 560 90 0 0 la_data_in[33]
port 198 nsew
flabel metal2 s 246366 -960 246478 480 0 FreeSans 560 90 0 0 la_data_in[34]
port 199 nsew
flabel metal2 s 249954 -960 250066 480 0 FreeSans 560 90 0 0 la_data_in[35]
port 200 nsew
flabel metal2 s 253450 -960 253562 480 0 FreeSans 560 90 0 0 la_data_in[36]
port 201 nsew
flabel metal2 s 257038 -960 257150 480 0 FreeSans 560 90 0 0 la_data_in[37]
port 202 nsew
flabel metal2 s 260626 -960 260738 480 0 FreeSans 560 90 0 0 la_data_in[38]
port 203 nsew
flabel metal2 s 264122 -960 264234 480 0 FreeSans 560 90 0 0 la_data_in[39]
port 204 nsew
flabel metal2 s 136426 -960 136538 480 0 FreeSans 560 90 0 0 la_data_in[3]
port 205 nsew
flabel metal2 s 267710 -960 267822 480 0 FreeSans 560 90 0 0 la_data_in[40]
port 206 nsew
flabel metal2 s 271206 -960 271318 480 0 FreeSans 560 90 0 0 la_data_in[41]
port 207 nsew
flabel metal2 s 274794 -960 274906 480 0 FreeSans 560 90 0 0 la_data_in[42]
port 208 nsew
flabel metal2 s 278290 -960 278402 480 0 FreeSans 560 90 0 0 la_data_in[43]
port 209 nsew
flabel metal2 s 281878 -960 281990 480 0 FreeSans 560 90 0 0 la_data_in[44]
port 210 nsew
flabel metal2 s 285374 -960 285486 480 0 FreeSans 560 90 0 0 la_data_in[45]
port 211 nsew
flabel metal2 s 288962 -960 289074 480 0 FreeSans 560 90 0 0 la_data_in[46]
port 212 nsew
flabel metal2 s 292550 -960 292662 480 0 FreeSans 560 90 0 0 la_data_in[47]
port 213 nsew
flabel metal2 s 296046 -960 296158 480 0 FreeSans 560 90 0 0 la_data_in[48]
port 214 nsew
flabel metal2 s 299634 -960 299746 480 0 FreeSans 560 90 0 0 la_data_in[49]
port 215 nsew
flabel metal2 s 140014 -960 140126 480 0 FreeSans 560 90 0 0 la_data_in[4]
port 216 nsew
flabel metal2 s 303130 -960 303242 480 0 FreeSans 560 90 0 0 la_data_in[50]
port 217 nsew
flabel metal2 s 306718 -960 306830 480 0 FreeSans 560 90 0 0 la_data_in[51]
port 218 nsew
flabel metal2 s 310214 -960 310326 480 0 FreeSans 560 90 0 0 la_data_in[52]
port 219 nsew
flabel metal2 s 313802 -960 313914 480 0 FreeSans 560 90 0 0 la_data_in[53]
port 220 nsew
flabel metal2 s 317298 -960 317410 480 0 FreeSans 560 90 0 0 la_data_in[54]
port 221 nsew
flabel metal2 s 320886 -960 320998 480 0 FreeSans 560 90 0 0 la_data_in[55]
port 222 nsew
flabel metal2 s 324382 -960 324494 480 0 FreeSans 560 90 0 0 la_data_in[56]
port 223 nsew
flabel metal2 s 327970 -960 328082 480 0 FreeSans 560 90 0 0 la_data_in[57]
port 224 nsew
flabel metal2 s 331558 -960 331670 480 0 FreeSans 560 90 0 0 la_data_in[58]
port 225 nsew
flabel metal2 s 335054 -960 335166 480 0 FreeSans 560 90 0 0 la_data_in[59]
port 226 nsew
flabel metal2 s 143510 -960 143622 480 0 FreeSans 560 90 0 0 la_data_in[5]
port 227 nsew
flabel metal2 s 338642 -960 338754 480 0 FreeSans 560 90 0 0 la_data_in[60]
port 228 nsew
flabel metal2 s 342138 -960 342250 480 0 FreeSans 560 90 0 0 la_data_in[61]
port 229 nsew
flabel metal2 s 345726 -960 345838 480 0 FreeSans 560 90 0 0 la_data_in[62]
port 230 nsew
flabel metal2 s 349222 -960 349334 480 0 FreeSans 560 90 0 0 la_data_in[63]
port 231 nsew
flabel metal2 s 352810 -960 352922 480 0 FreeSans 560 90 0 0 la_data_in[64]
port 232 nsew
flabel metal2 s 356306 -960 356418 480 0 FreeSans 560 90 0 0 la_data_in[65]
port 233 nsew
flabel metal2 s 359894 -960 360006 480 0 FreeSans 560 90 0 0 la_data_in[66]
port 234 nsew
flabel metal2 s 363482 -960 363594 480 0 FreeSans 560 90 0 0 la_data_in[67]
port 235 nsew
flabel metal2 s 366978 -960 367090 480 0 FreeSans 560 90 0 0 la_data_in[68]
port 236 nsew
flabel metal2 s 370566 -960 370678 480 0 FreeSans 560 90 0 0 la_data_in[69]
port 237 nsew
flabel metal2 s 147098 -960 147210 480 0 FreeSans 560 90 0 0 la_data_in[6]
port 238 nsew
flabel metal2 s 374062 -960 374174 480 0 FreeSans 560 90 0 0 la_data_in[70]
port 239 nsew
flabel metal2 s 377650 -960 377762 480 0 FreeSans 560 90 0 0 la_data_in[71]
port 240 nsew
flabel metal2 s 381146 -960 381258 480 0 FreeSans 560 90 0 0 la_data_in[72]
port 241 nsew
flabel metal2 s 384734 -960 384846 480 0 FreeSans 560 90 0 0 la_data_in[73]
port 242 nsew
flabel metal2 s 388230 -960 388342 480 0 FreeSans 560 90 0 0 la_data_in[74]
port 243 nsew
flabel metal2 s 391818 -960 391930 480 0 FreeSans 560 90 0 0 la_data_in[75]
port 244 nsew
flabel metal2 s 395314 -960 395426 480 0 FreeSans 560 90 0 0 la_data_in[76]
port 245 nsew
flabel metal2 s 398902 -960 399014 480 0 FreeSans 560 90 0 0 la_data_in[77]
port 246 nsew
flabel metal2 s 402490 -960 402602 480 0 FreeSans 560 90 0 0 la_data_in[78]
port 247 nsew
flabel metal2 s 405986 -960 406098 480 0 FreeSans 560 90 0 0 la_data_in[79]
port 248 nsew
flabel metal2 s 150594 -960 150706 480 0 FreeSans 560 90 0 0 la_data_in[7]
port 249 nsew
flabel metal2 s 409574 -960 409686 480 0 FreeSans 560 90 0 0 la_data_in[80]
port 250 nsew
flabel metal2 s 413070 -960 413182 480 0 FreeSans 560 90 0 0 la_data_in[81]
port 251 nsew
flabel metal2 s 416658 -960 416770 480 0 FreeSans 560 90 0 0 la_data_in[82]
port 252 nsew
flabel metal2 s 420154 -960 420266 480 0 FreeSans 560 90 0 0 la_data_in[83]
port 253 nsew
flabel metal2 s 423742 -960 423854 480 0 FreeSans 560 90 0 0 la_data_in[84]
port 254 nsew
flabel metal2 s 427238 -960 427350 480 0 FreeSans 560 90 0 0 la_data_in[85]
port 255 nsew
flabel metal2 s 430826 -960 430938 480 0 FreeSans 560 90 0 0 la_data_in[86]
port 256 nsew
flabel metal2 s 434414 -960 434526 480 0 FreeSans 560 90 0 0 la_data_in[87]
port 257 nsew
flabel metal2 s 437910 -960 438022 480 0 FreeSans 560 90 0 0 la_data_in[88]
port 258 nsew
flabel metal2 s 441498 -960 441610 480 0 FreeSans 560 90 0 0 la_data_in[89]
port 259 nsew
flabel metal2 s 154182 -960 154294 480 0 FreeSans 560 90 0 0 la_data_in[8]
port 260 nsew
flabel metal2 s 444994 -960 445106 480 0 FreeSans 560 90 0 0 la_data_in[90]
port 261 nsew
flabel metal2 s 448582 -960 448694 480 0 FreeSans 560 90 0 0 la_data_in[91]
port 262 nsew
flabel metal2 s 452078 -960 452190 480 0 FreeSans 560 90 0 0 la_data_in[92]
port 263 nsew
flabel metal2 s 455666 -960 455778 480 0 FreeSans 560 90 0 0 la_data_in[93]
port 264 nsew
flabel metal2 s 459162 -960 459274 480 0 FreeSans 560 90 0 0 la_data_in[94]
port 265 nsew
flabel metal2 s 462750 -960 462862 480 0 FreeSans 560 90 0 0 la_data_in[95]
port 266 nsew
flabel metal2 s 466246 -960 466358 480 0 FreeSans 560 90 0 0 la_data_in[96]
port 267 nsew
flabel metal2 s 469834 -960 469946 480 0 FreeSans 560 90 0 0 la_data_in[97]
port 268 nsew
flabel metal2 s 473422 -960 473534 480 0 FreeSans 560 90 0 0 la_data_in[98]
port 269 nsew
flabel metal2 s 476918 -960 477030 480 0 FreeSans 560 90 0 0 la_data_in[99]
port 270 nsew
flabel metal2 s 157770 -960 157882 480 0 FreeSans 560 90 0 0 la_data_in[9]
port 271 nsew
flabel metal2 s 126950 -960 127062 480 0 FreeSans 560 90 0 0 la_data_out[0]
port 272 nsew
flabel metal2 s 481702 -960 481814 480 0 FreeSans 560 90 0 0 la_data_out[100]
port 273 nsew
flabel metal2 s 485198 -960 485310 480 0 FreeSans 560 90 0 0 la_data_out[101]
port 274 nsew
flabel metal2 s 488786 -960 488898 480 0 FreeSans 560 90 0 0 la_data_out[102]
port 275 nsew
flabel metal2 s 492282 -960 492394 480 0 FreeSans 560 90 0 0 la_data_out[103]
port 276 nsew
flabel metal2 s 495870 -960 495982 480 0 FreeSans 560 90 0 0 la_data_out[104]
port 277 nsew
flabel metal2 s 499366 -960 499478 480 0 FreeSans 560 90 0 0 la_data_out[105]
port 278 nsew
flabel metal2 s 502954 -960 503066 480 0 FreeSans 560 90 0 0 la_data_out[106]
port 279 nsew
flabel metal2 s 506450 -960 506562 480 0 FreeSans 560 90 0 0 la_data_out[107]
port 280 nsew
flabel metal2 s 510038 -960 510150 480 0 FreeSans 560 90 0 0 la_data_out[108]
port 281 nsew
flabel metal2 s 513534 -960 513646 480 0 FreeSans 560 90 0 0 la_data_out[109]
port 282 nsew
flabel metal2 s 162462 -960 162574 480 0 FreeSans 560 90 0 0 la_data_out[10]
port 283 nsew
flabel metal2 s 517122 -960 517234 480 0 FreeSans 560 90 0 0 la_data_out[110]
port 284 nsew
flabel metal2 s 520710 -960 520822 480 0 FreeSans 560 90 0 0 la_data_out[111]
port 285 nsew
flabel metal2 s 524206 -960 524318 480 0 FreeSans 560 90 0 0 la_data_out[112]
port 286 nsew
flabel metal2 s 527794 -960 527906 480 0 FreeSans 560 90 0 0 la_data_out[113]
port 287 nsew
flabel metal2 s 531290 -960 531402 480 0 FreeSans 560 90 0 0 la_data_out[114]
port 288 nsew
flabel metal2 s 534878 -960 534990 480 0 FreeSans 560 90 0 0 la_data_out[115]
port 289 nsew
flabel metal2 s 538374 -960 538486 480 0 FreeSans 560 90 0 0 la_data_out[116]
port 290 nsew
flabel metal2 s 541962 -960 542074 480 0 FreeSans 560 90 0 0 la_data_out[117]
port 291 nsew
flabel metal2 s 545458 -960 545570 480 0 FreeSans 560 90 0 0 la_data_out[118]
port 292 nsew
flabel metal2 s 549046 -960 549158 480 0 FreeSans 560 90 0 0 la_data_out[119]
port 293 nsew
flabel metal2 s 166050 -960 166162 480 0 FreeSans 560 90 0 0 la_data_out[11]
port 294 nsew
flabel metal2 s 552634 -960 552746 480 0 FreeSans 560 90 0 0 la_data_out[120]
port 295 nsew
flabel metal2 s 556130 -960 556242 480 0 FreeSans 560 90 0 0 la_data_out[121]
port 296 nsew
flabel metal2 s 559718 -960 559830 480 0 FreeSans 560 90 0 0 la_data_out[122]
port 297 nsew
flabel metal2 s 563214 -960 563326 480 0 FreeSans 560 90 0 0 la_data_out[123]
port 298 nsew
flabel metal2 s 566802 -960 566914 480 0 FreeSans 560 90 0 0 la_data_out[124]
port 299 nsew
flabel metal2 s 570298 -960 570410 480 0 FreeSans 560 90 0 0 la_data_out[125]
port 300 nsew
flabel metal2 s 573886 -960 573998 480 0 FreeSans 560 90 0 0 la_data_out[126]
port 301 nsew
flabel metal2 s 577382 -960 577494 480 0 FreeSans 560 90 0 0 la_data_out[127]
port 302 nsew
flabel metal2 s 169546 -960 169658 480 0 FreeSans 560 90 0 0 la_data_out[12]
port 303 nsew
flabel metal2 s 173134 -960 173246 480 0 FreeSans 560 90 0 0 la_data_out[13]
port 304 nsew
flabel metal2 s 176630 -960 176742 480 0 FreeSans 560 90 0 0 la_data_out[14]
port 305 nsew
flabel metal2 s 180218 -960 180330 480 0 FreeSans 560 90 0 0 la_data_out[15]
port 306 nsew
flabel metal2 s 183714 -960 183826 480 0 FreeSans 560 90 0 0 la_data_out[16]
port 307 nsew
flabel metal2 s 187302 -960 187414 480 0 FreeSans 560 90 0 0 la_data_out[17]
port 308 nsew
flabel metal2 s 190798 -960 190910 480 0 FreeSans 560 90 0 0 la_data_out[18]
port 309 nsew
flabel metal2 s 194386 -960 194498 480 0 FreeSans 560 90 0 0 la_data_out[19]
port 310 nsew
flabel metal2 s 130538 -960 130650 480 0 FreeSans 560 90 0 0 la_data_out[1]
port 311 nsew
flabel metal2 s 197882 -960 197994 480 0 FreeSans 560 90 0 0 la_data_out[20]
port 312 nsew
flabel metal2 s 201470 -960 201582 480 0 FreeSans 560 90 0 0 la_data_out[21]
port 313 nsew
flabel metal2 s 205058 -960 205170 480 0 FreeSans 560 90 0 0 la_data_out[22]
port 314 nsew
flabel metal2 s 208554 -960 208666 480 0 FreeSans 560 90 0 0 la_data_out[23]
port 315 nsew
flabel metal2 s 212142 -960 212254 480 0 FreeSans 560 90 0 0 la_data_out[24]
port 316 nsew
flabel metal2 s 215638 -960 215750 480 0 FreeSans 560 90 0 0 la_data_out[25]
port 317 nsew
flabel metal2 s 219226 -960 219338 480 0 FreeSans 560 90 0 0 la_data_out[26]
port 318 nsew
flabel metal2 s 222722 -960 222834 480 0 FreeSans 560 90 0 0 la_data_out[27]
port 319 nsew
flabel metal2 s 226310 -960 226422 480 0 FreeSans 560 90 0 0 la_data_out[28]
port 320 nsew
flabel metal2 s 229806 -960 229918 480 0 FreeSans 560 90 0 0 la_data_out[29]
port 321 nsew
flabel metal2 s 134126 -960 134238 480 0 FreeSans 560 90 0 0 la_data_out[2]
port 322 nsew
flabel metal2 s 233394 -960 233506 480 0 FreeSans 560 90 0 0 la_data_out[30]
port 323 nsew
flabel metal2 s 236982 -960 237094 480 0 FreeSans 560 90 0 0 la_data_out[31]
port 324 nsew
flabel metal2 s 240478 -960 240590 480 0 FreeSans 560 90 0 0 la_data_out[32]
port 325 nsew
flabel metal2 s 244066 -960 244178 480 0 FreeSans 560 90 0 0 la_data_out[33]
port 326 nsew
flabel metal2 s 247562 -960 247674 480 0 FreeSans 560 90 0 0 la_data_out[34]
port 327 nsew
flabel metal2 s 251150 -960 251262 480 0 FreeSans 560 90 0 0 la_data_out[35]
port 328 nsew
flabel metal2 s 254646 -960 254758 480 0 FreeSans 560 90 0 0 la_data_out[36]
port 329 nsew
flabel metal2 s 258234 -960 258346 480 0 FreeSans 560 90 0 0 la_data_out[37]
port 330 nsew
flabel metal2 s 261730 -960 261842 480 0 FreeSans 560 90 0 0 la_data_out[38]
port 331 nsew
flabel metal2 s 265318 -960 265430 480 0 FreeSans 560 90 0 0 la_data_out[39]
port 332 nsew
flabel metal2 s 137622 -960 137734 480 0 FreeSans 560 90 0 0 la_data_out[3]
port 333 nsew
flabel metal2 s 268814 -960 268926 480 0 FreeSans 560 90 0 0 la_data_out[40]
port 334 nsew
flabel metal2 s 272402 -960 272514 480 0 FreeSans 560 90 0 0 la_data_out[41]
port 335 nsew
flabel metal2 s 275990 -960 276102 480 0 FreeSans 560 90 0 0 la_data_out[42]
port 336 nsew
flabel metal2 s 279486 -960 279598 480 0 FreeSans 560 90 0 0 la_data_out[43]
port 337 nsew
flabel metal2 s 283074 -960 283186 480 0 FreeSans 560 90 0 0 la_data_out[44]
port 338 nsew
flabel metal2 s 286570 -960 286682 480 0 FreeSans 560 90 0 0 la_data_out[45]
port 339 nsew
flabel metal2 s 290158 -960 290270 480 0 FreeSans 560 90 0 0 la_data_out[46]
port 340 nsew
flabel metal2 s 293654 -960 293766 480 0 FreeSans 560 90 0 0 la_data_out[47]
port 341 nsew
flabel metal2 s 297242 -960 297354 480 0 FreeSans 560 90 0 0 la_data_out[48]
port 342 nsew
flabel metal2 s 300738 -960 300850 480 0 FreeSans 560 90 0 0 la_data_out[49]
port 343 nsew
flabel metal2 s 141210 -960 141322 480 0 FreeSans 560 90 0 0 la_data_out[4]
port 344 nsew
flabel metal2 s 304326 -960 304438 480 0 FreeSans 560 90 0 0 la_data_out[50]
port 345 nsew
flabel metal2 s 307914 -960 308026 480 0 FreeSans 560 90 0 0 la_data_out[51]
port 346 nsew
flabel metal2 s 311410 -960 311522 480 0 FreeSans 560 90 0 0 la_data_out[52]
port 347 nsew
flabel metal2 s 314998 -960 315110 480 0 FreeSans 560 90 0 0 la_data_out[53]
port 348 nsew
flabel metal2 s 318494 -960 318606 480 0 FreeSans 560 90 0 0 la_data_out[54]
port 349 nsew
flabel metal2 s 322082 -960 322194 480 0 FreeSans 560 90 0 0 la_data_out[55]
port 350 nsew
flabel metal2 s 325578 -960 325690 480 0 FreeSans 560 90 0 0 la_data_out[56]
port 351 nsew
flabel metal2 s 329166 -960 329278 480 0 FreeSans 560 90 0 0 la_data_out[57]
port 352 nsew
flabel metal2 s 332662 -960 332774 480 0 FreeSans 560 90 0 0 la_data_out[58]
port 353 nsew
flabel metal2 s 336250 -960 336362 480 0 FreeSans 560 90 0 0 la_data_out[59]
port 354 nsew
flabel metal2 s 144706 -960 144818 480 0 FreeSans 560 90 0 0 la_data_out[5]
port 355 nsew
flabel metal2 s 339838 -960 339950 480 0 FreeSans 560 90 0 0 la_data_out[60]
port 356 nsew
flabel metal2 s 343334 -960 343446 480 0 FreeSans 560 90 0 0 la_data_out[61]
port 357 nsew
flabel metal2 s 346922 -960 347034 480 0 FreeSans 560 90 0 0 la_data_out[62]
port 358 nsew
flabel metal2 s 350418 -960 350530 480 0 FreeSans 560 90 0 0 la_data_out[63]
port 359 nsew
flabel metal2 s 354006 -960 354118 480 0 FreeSans 560 90 0 0 la_data_out[64]
port 360 nsew
flabel metal2 s 357502 -960 357614 480 0 FreeSans 560 90 0 0 la_data_out[65]
port 361 nsew
flabel metal2 s 361090 -960 361202 480 0 FreeSans 560 90 0 0 la_data_out[66]
port 362 nsew
flabel metal2 s 364586 -960 364698 480 0 FreeSans 560 90 0 0 la_data_out[67]
port 363 nsew
flabel metal2 s 368174 -960 368286 480 0 FreeSans 560 90 0 0 la_data_out[68]
port 364 nsew
flabel metal2 s 371670 -960 371782 480 0 FreeSans 560 90 0 0 la_data_out[69]
port 365 nsew
flabel metal2 s 148294 -960 148406 480 0 FreeSans 560 90 0 0 la_data_out[6]
port 366 nsew
flabel metal2 s 375258 -960 375370 480 0 FreeSans 560 90 0 0 la_data_out[70]
port 367 nsew
flabel metal2 s 378846 -960 378958 480 0 FreeSans 560 90 0 0 la_data_out[71]
port 368 nsew
flabel metal2 s 382342 -960 382454 480 0 FreeSans 560 90 0 0 la_data_out[72]
port 369 nsew
flabel metal2 s 385930 -960 386042 480 0 FreeSans 560 90 0 0 la_data_out[73]
port 370 nsew
flabel metal2 s 389426 -960 389538 480 0 FreeSans 560 90 0 0 la_data_out[74]
port 371 nsew
flabel metal2 s 393014 -960 393126 480 0 FreeSans 560 90 0 0 la_data_out[75]
port 372 nsew
flabel metal2 s 396510 -960 396622 480 0 FreeSans 560 90 0 0 la_data_out[76]
port 373 nsew
flabel metal2 s 400098 -960 400210 480 0 FreeSans 560 90 0 0 la_data_out[77]
port 374 nsew
flabel metal2 s 403594 -960 403706 480 0 FreeSans 560 90 0 0 la_data_out[78]
port 375 nsew
flabel metal2 s 407182 -960 407294 480 0 FreeSans 560 90 0 0 la_data_out[79]
port 376 nsew
flabel metal2 s 151790 -960 151902 480 0 FreeSans 560 90 0 0 la_data_out[7]
port 377 nsew
flabel metal2 s 410770 -960 410882 480 0 FreeSans 560 90 0 0 la_data_out[80]
port 378 nsew
flabel metal2 s 414266 -960 414378 480 0 FreeSans 560 90 0 0 la_data_out[81]
port 379 nsew
flabel metal2 s 417854 -960 417966 480 0 FreeSans 560 90 0 0 la_data_out[82]
port 380 nsew
flabel metal2 s 421350 -960 421462 480 0 FreeSans 560 90 0 0 la_data_out[83]
port 381 nsew
flabel metal2 s 424938 -960 425050 480 0 FreeSans 560 90 0 0 la_data_out[84]
port 382 nsew
flabel metal2 s 428434 -960 428546 480 0 FreeSans 560 90 0 0 la_data_out[85]
port 383 nsew
flabel metal2 s 432022 -960 432134 480 0 FreeSans 560 90 0 0 la_data_out[86]
port 384 nsew
flabel metal2 s 435518 -960 435630 480 0 FreeSans 560 90 0 0 la_data_out[87]
port 385 nsew
flabel metal2 s 439106 -960 439218 480 0 FreeSans 560 90 0 0 la_data_out[88]
port 386 nsew
flabel metal2 s 442602 -960 442714 480 0 FreeSans 560 90 0 0 la_data_out[89]
port 387 nsew
flabel metal2 s 155378 -960 155490 480 0 FreeSans 560 90 0 0 la_data_out[8]
port 388 nsew
flabel metal2 s 446190 -960 446302 480 0 FreeSans 560 90 0 0 la_data_out[90]
port 389 nsew
flabel metal2 s 449778 -960 449890 480 0 FreeSans 560 90 0 0 la_data_out[91]
port 390 nsew
flabel metal2 s 453274 -960 453386 480 0 FreeSans 560 90 0 0 la_data_out[92]
port 391 nsew
flabel metal2 s 456862 -960 456974 480 0 FreeSans 560 90 0 0 la_data_out[93]
port 392 nsew
flabel metal2 s 460358 -960 460470 480 0 FreeSans 560 90 0 0 la_data_out[94]
port 393 nsew
flabel metal2 s 463946 -960 464058 480 0 FreeSans 560 90 0 0 la_data_out[95]
port 394 nsew
flabel metal2 s 467442 -960 467554 480 0 FreeSans 560 90 0 0 la_data_out[96]
port 395 nsew
flabel metal2 s 471030 -960 471142 480 0 FreeSans 560 90 0 0 la_data_out[97]
port 396 nsew
flabel metal2 s 474526 -960 474638 480 0 FreeSans 560 90 0 0 la_data_out[98]
port 397 nsew
flabel metal2 s 478114 -960 478226 480 0 FreeSans 560 90 0 0 la_data_out[99]
port 398 nsew
flabel metal2 s 158874 -960 158986 480 0 FreeSans 560 90 0 0 la_data_out[9]
port 399 nsew
flabel metal2 s 128146 -960 128258 480 0 FreeSans 560 90 0 0 la_oenb[0]
port 400 nsew
flabel metal2 s 482806 -960 482918 480 0 FreeSans 560 90 0 0 la_oenb[100]
port 401 nsew
flabel metal2 s 486394 -960 486506 480 0 FreeSans 560 90 0 0 la_oenb[101]
port 402 nsew
flabel metal2 s 489890 -960 490002 480 0 FreeSans 560 90 0 0 la_oenb[102]
port 403 nsew
flabel metal2 s 493478 -960 493590 480 0 FreeSans 560 90 0 0 la_oenb[103]
port 404 nsew
flabel metal2 s 497066 -960 497178 480 0 FreeSans 560 90 0 0 la_oenb[104]
port 405 nsew
flabel metal2 s 500562 -960 500674 480 0 FreeSans 560 90 0 0 la_oenb[105]
port 406 nsew
flabel metal2 s 504150 -960 504262 480 0 FreeSans 560 90 0 0 la_oenb[106]
port 407 nsew
flabel metal2 s 507646 -960 507758 480 0 FreeSans 560 90 0 0 la_oenb[107]
port 408 nsew
flabel metal2 s 511234 -960 511346 480 0 FreeSans 560 90 0 0 la_oenb[108]
port 409 nsew
flabel metal2 s 514730 -960 514842 480 0 FreeSans 560 90 0 0 la_oenb[109]
port 410 nsew
flabel metal2 s 163658 -960 163770 480 0 FreeSans 560 90 0 0 la_oenb[10]
port 411 nsew
flabel metal2 s 518318 -960 518430 480 0 FreeSans 560 90 0 0 la_oenb[110]
port 412 nsew
flabel metal2 s 521814 -960 521926 480 0 FreeSans 560 90 0 0 la_oenb[111]
port 413 nsew
flabel metal2 s 525402 -960 525514 480 0 FreeSans 560 90 0 0 la_oenb[112]
port 414 nsew
flabel metal2 s 528990 -960 529102 480 0 FreeSans 560 90 0 0 la_oenb[113]
port 415 nsew
flabel metal2 s 532486 -960 532598 480 0 FreeSans 560 90 0 0 la_oenb[114]
port 416 nsew
flabel metal2 s 536074 -960 536186 480 0 FreeSans 560 90 0 0 la_oenb[115]
port 417 nsew
flabel metal2 s 539570 -960 539682 480 0 FreeSans 560 90 0 0 la_oenb[116]
port 418 nsew
flabel metal2 s 543158 -960 543270 480 0 FreeSans 560 90 0 0 la_oenb[117]
port 419 nsew
flabel metal2 s 546654 -960 546766 480 0 FreeSans 560 90 0 0 la_oenb[118]
port 420 nsew
flabel metal2 s 550242 -960 550354 480 0 FreeSans 560 90 0 0 la_oenb[119]
port 421 nsew
flabel metal2 s 167154 -960 167266 480 0 FreeSans 560 90 0 0 la_oenb[11]
port 422 nsew
flabel metal2 s 553738 -960 553850 480 0 FreeSans 560 90 0 0 la_oenb[120]
port 423 nsew
flabel metal2 s 557326 -960 557438 480 0 FreeSans 560 90 0 0 la_oenb[121]
port 424 nsew
flabel metal2 s 560822 -960 560934 480 0 FreeSans 560 90 0 0 la_oenb[122]
port 425 nsew
flabel metal2 s 564410 -960 564522 480 0 FreeSans 560 90 0 0 la_oenb[123]
port 426 nsew
flabel metal2 s 567998 -960 568110 480 0 FreeSans 560 90 0 0 la_oenb[124]
port 427 nsew
flabel metal2 s 571494 -960 571606 480 0 FreeSans 560 90 0 0 la_oenb[125]
port 428 nsew
flabel metal2 s 575082 -960 575194 480 0 FreeSans 560 90 0 0 la_oenb[126]
port 429 nsew
flabel metal2 s 578578 -960 578690 480 0 FreeSans 560 90 0 0 la_oenb[127]
port 430 nsew
flabel metal2 s 170742 -960 170854 480 0 FreeSans 560 90 0 0 la_oenb[12]
port 431 nsew
flabel metal2 s 174238 -960 174350 480 0 FreeSans 560 90 0 0 la_oenb[13]
port 432 nsew
flabel metal2 s 177826 -960 177938 480 0 FreeSans 560 90 0 0 la_oenb[14]
port 433 nsew
flabel metal2 s 181414 -960 181526 480 0 FreeSans 560 90 0 0 la_oenb[15]
port 434 nsew
flabel metal2 s 184910 -960 185022 480 0 FreeSans 560 90 0 0 la_oenb[16]
port 435 nsew
flabel metal2 s 188498 -960 188610 480 0 FreeSans 560 90 0 0 la_oenb[17]
port 436 nsew
flabel metal2 s 191994 -960 192106 480 0 FreeSans 560 90 0 0 la_oenb[18]
port 437 nsew
flabel metal2 s 195582 -960 195694 480 0 FreeSans 560 90 0 0 la_oenb[19]
port 438 nsew
flabel metal2 s 131734 -960 131846 480 0 FreeSans 560 90 0 0 la_oenb[1]
port 439 nsew
flabel metal2 s 199078 -960 199190 480 0 FreeSans 560 90 0 0 la_oenb[20]
port 440 nsew
flabel metal2 s 202666 -960 202778 480 0 FreeSans 560 90 0 0 la_oenb[21]
port 441 nsew
flabel metal2 s 206162 -960 206274 480 0 FreeSans 560 90 0 0 la_oenb[22]
port 442 nsew
flabel metal2 s 209750 -960 209862 480 0 FreeSans 560 90 0 0 la_oenb[23]
port 443 nsew
flabel metal2 s 213338 -960 213450 480 0 FreeSans 560 90 0 0 la_oenb[24]
port 444 nsew
flabel metal2 s 216834 -960 216946 480 0 FreeSans 560 90 0 0 la_oenb[25]
port 445 nsew
flabel metal2 s 220422 -960 220534 480 0 FreeSans 560 90 0 0 la_oenb[26]
port 446 nsew
flabel metal2 s 223918 -960 224030 480 0 FreeSans 560 90 0 0 la_oenb[27]
port 447 nsew
flabel metal2 s 227506 -960 227618 480 0 FreeSans 560 90 0 0 la_oenb[28]
port 448 nsew
flabel metal2 s 231002 -960 231114 480 0 FreeSans 560 90 0 0 la_oenb[29]
port 449 nsew
flabel metal2 s 135230 -960 135342 480 0 FreeSans 560 90 0 0 la_oenb[2]
port 450 nsew
flabel metal2 s 234590 -960 234702 480 0 FreeSans 560 90 0 0 la_oenb[30]
port 451 nsew
flabel metal2 s 238086 -960 238198 480 0 FreeSans 560 90 0 0 la_oenb[31]
port 452 nsew
flabel metal2 s 241674 -960 241786 480 0 FreeSans 560 90 0 0 la_oenb[32]
port 453 nsew
flabel metal2 s 245170 -960 245282 480 0 FreeSans 560 90 0 0 la_oenb[33]
port 454 nsew
flabel metal2 s 248758 -960 248870 480 0 FreeSans 560 90 0 0 la_oenb[34]
port 455 nsew
flabel metal2 s 252346 -960 252458 480 0 FreeSans 560 90 0 0 la_oenb[35]
port 456 nsew
flabel metal2 s 255842 -960 255954 480 0 FreeSans 560 90 0 0 la_oenb[36]
port 457 nsew
flabel metal2 s 259430 -960 259542 480 0 FreeSans 560 90 0 0 la_oenb[37]
port 458 nsew
flabel metal2 s 262926 -960 263038 480 0 FreeSans 560 90 0 0 la_oenb[38]
port 459 nsew
flabel metal2 s 266514 -960 266626 480 0 FreeSans 560 90 0 0 la_oenb[39]
port 460 nsew
flabel metal2 s 138818 -960 138930 480 0 FreeSans 560 90 0 0 la_oenb[3]
port 461 nsew
flabel metal2 s 270010 -960 270122 480 0 FreeSans 560 90 0 0 la_oenb[40]
port 462 nsew
flabel metal2 s 273598 -960 273710 480 0 FreeSans 560 90 0 0 la_oenb[41]
port 463 nsew
flabel metal2 s 277094 -960 277206 480 0 FreeSans 560 90 0 0 la_oenb[42]
port 464 nsew
flabel metal2 s 280682 -960 280794 480 0 FreeSans 560 90 0 0 la_oenb[43]
port 465 nsew
flabel metal2 s 284270 -960 284382 480 0 FreeSans 560 90 0 0 la_oenb[44]
port 466 nsew
flabel metal2 s 287766 -960 287878 480 0 FreeSans 560 90 0 0 la_oenb[45]
port 467 nsew
flabel metal2 s 291354 -960 291466 480 0 FreeSans 560 90 0 0 la_oenb[46]
port 468 nsew
flabel metal2 s 294850 -960 294962 480 0 FreeSans 560 90 0 0 la_oenb[47]
port 469 nsew
flabel metal2 s 298438 -960 298550 480 0 FreeSans 560 90 0 0 la_oenb[48]
port 470 nsew
flabel metal2 s 301934 -960 302046 480 0 FreeSans 560 90 0 0 la_oenb[49]
port 471 nsew
flabel metal2 s 142406 -960 142518 480 0 FreeSans 560 90 0 0 la_oenb[4]
port 472 nsew
flabel metal2 s 305522 -960 305634 480 0 FreeSans 560 90 0 0 la_oenb[50]
port 473 nsew
flabel metal2 s 309018 -960 309130 480 0 FreeSans 560 90 0 0 la_oenb[51]
port 474 nsew
flabel metal2 s 312606 -960 312718 480 0 FreeSans 560 90 0 0 la_oenb[52]
port 475 nsew
flabel metal2 s 316194 -960 316306 480 0 FreeSans 560 90 0 0 la_oenb[53]
port 476 nsew
flabel metal2 s 319690 -960 319802 480 0 FreeSans 560 90 0 0 la_oenb[54]
port 477 nsew
flabel metal2 s 323278 -960 323390 480 0 FreeSans 560 90 0 0 la_oenb[55]
port 478 nsew
flabel metal2 s 326774 -960 326886 480 0 FreeSans 560 90 0 0 la_oenb[56]
port 479 nsew
flabel metal2 s 330362 -960 330474 480 0 FreeSans 560 90 0 0 la_oenb[57]
port 480 nsew
flabel metal2 s 333858 -960 333970 480 0 FreeSans 560 90 0 0 la_oenb[58]
port 481 nsew
flabel metal2 s 337446 -960 337558 480 0 FreeSans 560 90 0 0 la_oenb[59]
port 482 nsew
flabel metal2 s 145902 -960 146014 480 0 FreeSans 560 90 0 0 la_oenb[5]
port 483 nsew
flabel metal2 s 340942 -960 341054 480 0 FreeSans 560 90 0 0 la_oenb[60]
port 484 nsew
flabel metal2 s 344530 -960 344642 480 0 FreeSans 560 90 0 0 la_oenb[61]
port 485 nsew
flabel metal2 s 348026 -960 348138 480 0 FreeSans 560 90 0 0 la_oenb[62]
port 486 nsew
flabel metal2 s 351614 -960 351726 480 0 FreeSans 560 90 0 0 la_oenb[63]
port 487 nsew
flabel metal2 s 355202 -960 355314 480 0 FreeSans 560 90 0 0 la_oenb[64]
port 488 nsew
flabel metal2 s 358698 -960 358810 480 0 FreeSans 560 90 0 0 la_oenb[65]
port 489 nsew
flabel metal2 s 362286 -960 362398 480 0 FreeSans 560 90 0 0 la_oenb[66]
port 490 nsew
flabel metal2 s 365782 -960 365894 480 0 FreeSans 560 90 0 0 la_oenb[67]
port 491 nsew
flabel metal2 s 369370 -960 369482 480 0 FreeSans 560 90 0 0 la_oenb[68]
port 492 nsew
flabel metal2 s 372866 -960 372978 480 0 FreeSans 560 90 0 0 la_oenb[69]
port 493 nsew
flabel metal2 s 149490 -960 149602 480 0 FreeSans 560 90 0 0 la_oenb[6]
port 494 nsew
flabel metal2 s 376454 -960 376566 480 0 FreeSans 560 90 0 0 la_oenb[70]
port 495 nsew
flabel metal2 s 379950 -960 380062 480 0 FreeSans 560 90 0 0 la_oenb[71]
port 496 nsew
flabel metal2 s 383538 -960 383650 480 0 FreeSans 560 90 0 0 la_oenb[72]
port 497 nsew
flabel metal2 s 387126 -960 387238 480 0 FreeSans 560 90 0 0 la_oenb[73]
port 498 nsew
flabel metal2 s 390622 -960 390734 480 0 FreeSans 560 90 0 0 la_oenb[74]
port 499 nsew
flabel metal2 s 394210 -960 394322 480 0 FreeSans 560 90 0 0 la_oenb[75]
port 500 nsew
flabel metal2 s 397706 -960 397818 480 0 FreeSans 560 90 0 0 la_oenb[76]
port 501 nsew
flabel metal2 s 401294 -960 401406 480 0 FreeSans 560 90 0 0 la_oenb[77]
port 502 nsew
flabel metal2 s 404790 -960 404902 480 0 FreeSans 560 90 0 0 la_oenb[78]
port 503 nsew
flabel metal2 s 408378 -960 408490 480 0 FreeSans 560 90 0 0 la_oenb[79]
port 504 nsew
flabel metal2 s 152986 -960 153098 480 0 FreeSans 560 90 0 0 la_oenb[7]
port 505 nsew
flabel metal2 s 411874 -960 411986 480 0 FreeSans 560 90 0 0 la_oenb[80]
port 506 nsew
flabel metal2 s 415462 -960 415574 480 0 FreeSans 560 90 0 0 la_oenb[81]
port 507 nsew
flabel metal2 s 418958 -960 419070 480 0 FreeSans 560 90 0 0 la_oenb[82]
port 508 nsew
flabel metal2 s 422546 -960 422658 480 0 FreeSans 560 90 0 0 la_oenb[83]
port 509 nsew
flabel metal2 s 426134 -960 426246 480 0 FreeSans 560 90 0 0 la_oenb[84]
port 510 nsew
flabel metal2 s 429630 -960 429742 480 0 FreeSans 560 90 0 0 la_oenb[85]
port 511 nsew
flabel metal2 s 433218 -960 433330 480 0 FreeSans 560 90 0 0 la_oenb[86]
port 512 nsew
flabel metal2 s 436714 -960 436826 480 0 FreeSans 560 90 0 0 la_oenb[87]
port 513 nsew
flabel metal2 s 440302 -960 440414 480 0 FreeSans 560 90 0 0 la_oenb[88]
port 514 nsew
flabel metal2 s 443798 -960 443910 480 0 FreeSans 560 90 0 0 la_oenb[89]
port 515 nsew
flabel metal2 s 156574 -960 156686 480 0 FreeSans 560 90 0 0 la_oenb[8]
port 516 nsew
flabel metal2 s 447386 -960 447498 480 0 FreeSans 560 90 0 0 la_oenb[90]
port 517 nsew
flabel metal2 s 450882 -960 450994 480 0 FreeSans 560 90 0 0 la_oenb[91]
port 518 nsew
flabel metal2 s 454470 -960 454582 480 0 FreeSans 560 90 0 0 la_oenb[92]
port 519 nsew
flabel metal2 s 458058 -960 458170 480 0 FreeSans 560 90 0 0 la_oenb[93]
port 520 nsew
flabel metal2 s 461554 -960 461666 480 0 FreeSans 560 90 0 0 la_oenb[94]
port 521 nsew
flabel metal2 s 465142 -960 465254 480 0 FreeSans 560 90 0 0 la_oenb[95]
port 522 nsew
flabel metal2 s 468638 -960 468750 480 0 FreeSans 560 90 0 0 la_oenb[96]
port 523 nsew
flabel metal2 s 472226 -960 472338 480 0 FreeSans 560 90 0 0 la_oenb[97]
port 524 nsew
flabel metal2 s 475722 -960 475834 480 0 FreeSans 560 90 0 0 la_oenb[98]
port 525 nsew
flabel metal2 s 479310 -960 479422 480 0 FreeSans 560 90 0 0 la_oenb[99]
port 526 nsew
flabel metal2 s 160070 -960 160182 480 0 FreeSans 560 90 0 0 la_oenb[9]
port 527 nsew
flabel metal2 s 579774 -960 579886 480 0 FreeSans 560 90 0 0 user_clock2
port 528 nsew
flabel metal2 s 580970 -960 581082 480 0 FreeSans 560 90 0 0 user_irq[0]
port 529 nsew
flabel metal2 s 582166 -960 582278 480 0 FreeSans 560 90 0 0 user_irq[1]
port 530 nsew
flabel metal2 s 583362 -960 583474 480 0 FreeSans 560 90 0 0 user_irq[2]
port 531 nsew
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 397794 -7654 398414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 361794 -7654 362414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 325794 -7654 326414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 289794 -7654 290414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 253794 282628 254414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 253794 -7654 254414 2988 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 217794 -7654 218414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 181794 -7654 182414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 145794 -7654 146414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 109794 -7654 110414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 73794 -7654 74414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 694306 592650 694926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 658306 592650 658926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 622306 592650 622926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 586306 592650 586926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 550306 592650 550926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 514306 592650 514926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 478306 592650 478926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 442306 592650 442926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 406306 592650 406926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 370306 592650 370926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 334306 592650 334926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 298306 592650 298926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 262306 592650 262926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 226306 592650 226926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 190306 592650 190926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 154306 592650 154926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 118306 592650 118926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 82306 592650 82926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 46306 592650 46926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 10306 592650 10926 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal4 s 549234 -7654 549854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 513234 -7654 513854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 477234 -7654 477854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 441234 -7654 441854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 405234 -7654 405854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 369234 -7654 369854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 333234 -7654 333854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 297234 -7654 297854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 261234 282628 261854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 261234 -7654 261854 2988 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 225234 -7654 225854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 189234 -7654 189854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 153234 -7654 153854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 117234 -7654 117854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 81234 -7654 81854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 45234 -7654 45854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 9234 -7654 9854 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 665746 592650 666366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 629746 592650 630366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 593746 592650 594366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 557746 592650 558366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 521746 592650 522366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 485746 592650 486366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 449746 592650 450366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 413746 592650 414366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 377746 592650 378366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 341746 592650 342366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 305746 592650 306366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 269746 592650 270366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 233746 592650 234366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 197746 592650 198366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 161746 592650 162366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 125746 592650 126366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 89746 592650 90366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 53746 592650 54366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 17746 592650 18366 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal4 s 556674 -7654 557294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 520674 -7654 521294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 484674 -7654 485294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 448674 -7654 449294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 412674 -7654 413294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 376674 -7654 377294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 340674 -7654 341294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 304674 -7654 305294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 268674 -7654 269294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 232674 -7654 233294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 196674 -7654 197294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 160674 -7654 161294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 124674 -7654 125294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 88674 -7654 89294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 52674 -7654 53294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 16674 149892 17294 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 16674 -7654 17294 4076 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 673186 592650 673806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 637186 592650 637806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 601186 592650 601806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 565186 592650 565806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 529186 592650 529806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 493186 592650 493806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 457186 592650 457806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 421186 592650 421806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 385186 592650 385806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 349186 592650 349806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 313186 592650 313806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 277186 592650 277806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 241186 592650 241806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 205186 592650 205806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 169186 592650 169806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 133186 592650 133806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 97186 592650 97806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 61186 592650 61806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 25186 592650 25806 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal4 s 564114 -7654 564734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 528114 -7654 528734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 492114 -7654 492734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 456114 -7654 456734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 420114 -7654 420734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 384114 -7654 384734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 348114 -7654 348734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 312114 -7654 312734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 276114 -7654 276734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 240114 -7654 240734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 204114 -7654 204734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 168114 -7654 168734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 132114 -7654 132734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 96114 -7654 96734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 60114 -7654 60734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 24114 282628 24734 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 24114 -7654 24734 2988 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 669466 592650 670086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 633466 592650 634086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 597466 592650 598086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 561466 592650 562086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 525466 592650 526086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 489466 592650 490086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 453466 592650 454086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 417466 592650 418086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 381466 592650 382086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 345466 592650 346086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 309466 592650 310086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 273466 592650 274086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 237466 592650 238086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 201466 592650 202086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 165466 592650 166086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 129466 592650 130086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 93466 592650 94086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 57466 592650 58086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 21466 592650 22086 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal4 s 560394 -7654 561014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 524394 -7654 525014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 488394 -7654 489014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 452394 -7654 453014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 416394 -7654 417014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 380394 -7654 381014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 344394 -7654 345014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 308394 -7654 309014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 272394 -7654 273014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 236394 -7654 237014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 200394 282628 201014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 200394 -7654 201014 2988 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 164394 -7654 165014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 128394 -7654 129014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 92394 282628 93014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 92394 -7654 93014 2988 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 56394 -7654 57014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 20394 -7654 21014 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 676906 592650 677526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 640906 592650 641526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 604906 592650 605526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 568906 592650 569526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 532906 592650 533526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 496906 592650 497526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 460906 592650 461526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 424906 592650 425526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 388906 592650 389526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 352906 592650 353526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 316906 592650 317526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 280906 592650 281526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 244906 592650 245526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 208906 592650 209526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 172906 592650 173526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 136906 592650 137526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 100906 592650 101526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 64906 592650 65526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 28906 592650 29526 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal4 s 567834 -7654 568454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 531834 -7654 532454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 495834 -7654 496454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 459834 -7654 460454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 423834 -7654 424454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 387834 -7654 388454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 351834 -7654 352454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 315834 -7654 316454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 279834 -7654 280454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 243834 -7654 244454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 207834 282628 208454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 207834 -7654 208454 2988 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 171834 -7654 172454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 135834 -7654 136454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 99834 -7654 100454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 63834 -7654 64454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 27834 -7654 28454 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 690586 592650 691206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 654586 592650 655206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 618586 592650 619206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 582586 592650 583206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 546586 592650 547206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 510586 592650 511206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 474586 592650 475206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 438586 592650 439206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 402586 592650 403206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 366586 592650 367206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 330586 592650 331206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 294586 592650 295206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 258586 592650 259206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 222586 592650 223206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 186586 592650 187206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 150586 592650 151206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 114586 592650 115206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 78586 592650 79206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 42586 592650 43206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 6586 592650 7206 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal4 s 581514 -7654 582134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 545514 -7654 546134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 509514 -7654 510134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 473514 -7654 474134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 437514 -7654 438134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 401514 -7654 402134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 365514 -7654 366134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 329514 -7654 330134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 293514 -7654 294134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 257514 -7654 258134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 221514 -7654 222134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 185514 282628 186134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 185514 -7654 186134 2988 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 149514 -7654 150134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 113514 146817 114134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 113514 -7654 114134 3207 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 77514 282628 78134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 77514 -7654 78134 2988 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 41514 -7654 42134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 5514 -7654 6134 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 698026 592650 698646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 662026 592650 662646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 626026 592650 626646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 590026 592650 590646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 554026 592650 554646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 518026 592650 518646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 482026 592650 482646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 446026 592650 446646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 410026 592650 410646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 374026 592650 374646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 338026 592650 338646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 302026 592650 302646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 266026 592650 266646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 230026 592650 230646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 194026 592650 194646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 158026 592650 158646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 122026 592650 122646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 86026 592650 86646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 50026 592650 50646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 14026 592650 14646 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal4 s 552954 -7654 553574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 516954 -7654 517574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 480954 -7654 481574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 444954 -7654 445574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 408954 -7654 409574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 372954 -7654 373574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 336954 -7654 337574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 300954 -7654 301574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 264954 -7654 265574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 228954 -7654 229574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 192954 282628 193574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 192954 -7654 193574 2988 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 156954 -7654 157574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 120954 -7654 121574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 84954 282628 85574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 84954 -7654 85574 2988 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 48954 -7654 49574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 12954 -7654 13574 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal2 s 542 -960 654 480 0 FreeSans 560 90 0 0 wb_clk_i
port 540 nsew
flabel metal2 s 1646 -960 1758 480 0 FreeSans 560 90 0 0 wb_rst_i
port 541 nsew
flabel metal2 s 2842 -960 2954 480 0 FreeSans 560 90 0 0 wbs_ack_o
port 542 nsew
flabel metal2 s 7626 -960 7738 480 0 FreeSans 560 90 0 0 wbs_adr_i[0]
port 543 nsew
flabel metal2 s 47830 -960 47942 480 0 FreeSans 560 90 0 0 wbs_adr_i[10]
port 544 nsew
flabel metal2 s 51326 -960 51438 480 0 FreeSans 560 90 0 0 wbs_adr_i[11]
port 545 nsew
flabel metal2 s 54914 -960 55026 480 0 FreeSans 560 90 0 0 wbs_adr_i[12]
port 546 nsew
flabel metal2 s 58410 -960 58522 480 0 FreeSans 560 90 0 0 wbs_adr_i[13]
port 547 nsew
flabel metal2 s 61998 -960 62110 480 0 FreeSans 560 90 0 0 wbs_adr_i[14]
port 548 nsew
flabel metal2 s 65494 -960 65606 480 0 FreeSans 560 90 0 0 wbs_adr_i[15]
port 549 nsew
flabel metal2 s 69082 -960 69194 480 0 FreeSans 560 90 0 0 wbs_adr_i[16]
port 550 nsew
flabel metal2 s 72578 -960 72690 480 0 FreeSans 560 90 0 0 wbs_adr_i[17]
port 551 nsew
flabel metal2 s 76166 -960 76278 480 0 FreeSans 560 90 0 0 wbs_adr_i[18]
port 552 nsew
flabel metal2 s 79662 -960 79774 480 0 FreeSans 560 90 0 0 wbs_adr_i[19]
port 553 nsew
flabel metal2 s 12318 -960 12430 480 0 FreeSans 560 90 0 0 wbs_adr_i[1]
port 554 nsew
flabel metal2 s 83250 -960 83362 480 0 FreeSans 560 90 0 0 wbs_adr_i[20]
port 555 nsew
flabel metal2 s 86838 -960 86950 480 0 FreeSans 560 90 0 0 wbs_adr_i[21]
port 556 nsew
flabel metal2 s 90334 -960 90446 480 0 FreeSans 560 90 0 0 wbs_adr_i[22]
port 557 nsew
flabel metal2 s 93922 -960 94034 480 0 FreeSans 560 90 0 0 wbs_adr_i[23]
port 558 nsew
flabel metal2 s 97418 -960 97530 480 0 FreeSans 560 90 0 0 wbs_adr_i[24]
port 559 nsew
flabel metal2 s 101006 -960 101118 480 0 FreeSans 560 90 0 0 wbs_adr_i[25]
port 560 nsew
flabel metal2 s 104502 -960 104614 480 0 FreeSans 560 90 0 0 wbs_adr_i[26]
port 561 nsew
flabel metal2 s 108090 -960 108202 480 0 FreeSans 560 90 0 0 wbs_adr_i[27]
port 562 nsew
flabel metal2 s 111586 -960 111698 480 0 FreeSans 560 90 0 0 wbs_adr_i[28]
port 563 nsew
flabel metal2 s 115174 -960 115286 480 0 FreeSans 560 90 0 0 wbs_adr_i[29]
port 564 nsew
flabel metal2 s 17010 -960 17122 480 0 FreeSans 560 90 0 0 wbs_adr_i[2]
port 565 nsew
flabel metal2 s 118762 -960 118874 480 0 FreeSans 560 90 0 0 wbs_adr_i[30]
port 566 nsew
flabel metal2 s 122258 -960 122370 480 0 FreeSans 560 90 0 0 wbs_adr_i[31]
port 567 nsew
flabel metal2 s 21794 -960 21906 480 0 FreeSans 560 90 0 0 wbs_adr_i[3]
port 568 nsew
flabel metal2 s 26486 -960 26598 480 0 FreeSans 560 90 0 0 wbs_adr_i[4]
port 569 nsew
flabel metal2 s 30074 -960 30186 480 0 FreeSans 560 90 0 0 wbs_adr_i[5]
port 570 nsew
flabel metal2 s 33570 -960 33682 480 0 FreeSans 560 90 0 0 wbs_adr_i[6]
port 571 nsew
flabel metal2 s 37158 -960 37270 480 0 FreeSans 560 90 0 0 wbs_adr_i[7]
port 572 nsew
flabel metal2 s 40654 -960 40766 480 0 FreeSans 560 90 0 0 wbs_adr_i[8]
port 573 nsew
flabel metal2 s 44242 -960 44354 480 0 FreeSans 560 90 0 0 wbs_adr_i[9]
port 574 nsew
flabel metal2 s 4038 -960 4150 480 0 FreeSans 560 90 0 0 wbs_cyc_i
port 575 nsew
flabel metal2 s 8730 -960 8842 480 0 FreeSans 560 90 0 0 wbs_dat_i[0]
port 576 nsew
flabel metal2 s 48934 -960 49046 480 0 FreeSans 560 90 0 0 wbs_dat_i[10]
port 577 nsew
flabel metal2 s 52522 -960 52634 480 0 FreeSans 560 90 0 0 wbs_dat_i[11]
port 578 nsew
flabel metal2 s 56018 -960 56130 480 0 FreeSans 560 90 0 0 wbs_dat_i[12]
port 579 nsew
flabel metal2 s 59606 -960 59718 480 0 FreeSans 560 90 0 0 wbs_dat_i[13]
port 580 nsew
flabel metal2 s 63194 -960 63306 480 0 FreeSans 560 90 0 0 wbs_dat_i[14]
port 581 nsew
flabel metal2 s 66690 -960 66802 480 0 FreeSans 560 90 0 0 wbs_dat_i[15]
port 582 nsew
flabel metal2 s 70278 -960 70390 480 0 FreeSans 560 90 0 0 wbs_dat_i[16]
port 583 nsew
flabel metal2 s 73774 -960 73886 480 0 FreeSans 560 90 0 0 wbs_dat_i[17]
port 584 nsew
flabel metal2 s 77362 -960 77474 480 0 FreeSans 560 90 0 0 wbs_dat_i[18]
port 585 nsew
flabel metal2 s 80858 -960 80970 480 0 FreeSans 560 90 0 0 wbs_dat_i[19]
port 586 nsew
flabel metal2 s 13514 -960 13626 480 0 FreeSans 560 90 0 0 wbs_dat_i[1]
port 587 nsew
flabel metal2 s 84446 -960 84558 480 0 FreeSans 560 90 0 0 wbs_dat_i[20]
port 588 nsew
flabel metal2 s 87942 -960 88054 480 0 FreeSans 560 90 0 0 wbs_dat_i[21]
port 589 nsew
flabel metal2 s 91530 -960 91642 480 0 FreeSans 560 90 0 0 wbs_dat_i[22]
port 590 nsew
flabel metal2 s 95118 -960 95230 480 0 FreeSans 560 90 0 0 wbs_dat_i[23]
port 591 nsew
flabel metal2 s 98614 -960 98726 480 0 FreeSans 560 90 0 0 wbs_dat_i[24]
port 592 nsew
flabel metal2 s 102202 -960 102314 480 0 FreeSans 560 90 0 0 wbs_dat_i[25]
port 593 nsew
flabel metal2 s 105698 -960 105810 480 0 FreeSans 560 90 0 0 wbs_dat_i[26]
port 594 nsew
flabel metal2 s 109286 -960 109398 480 0 FreeSans 560 90 0 0 wbs_dat_i[27]
port 595 nsew
flabel metal2 s 112782 -960 112894 480 0 FreeSans 560 90 0 0 wbs_dat_i[28]
port 596 nsew
flabel metal2 s 116370 -960 116482 480 0 FreeSans 560 90 0 0 wbs_dat_i[29]
port 597 nsew
flabel metal2 s 18206 -960 18318 480 0 FreeSans 560 90 0 0 wbs_dat_i[2]
port 598 nsew
flabel metal2 s 119866 -960 119978 480 0 FreeSans 560 90 0 0 wbs_dat_i[30]
port 599 nsew
flabel metal2 s 123454 -960 123566 480 0 FreeSans 560 90 0 0 wbs_dat_i[31]
port 600 nsew
flabel metal2 s 22990 -960 23102 480 0 FreeSans 560 90 0 0 wbs_dat_i[3]
port 601 nsew
flabel metal2 s 27682 -960 27794 480 0 FreeSans 560 90 0 0 wbs_dat_i[4]
port 602 nsew
flabel metal2 s 31270 -960 31382 480 0 FreeSans 560 90 0 0 wbs_dat_i[5]
port 603 nsew
flabel metal2 s 34766 -960 34878 480 0 FreeSans 560 90 0 0 wbs_dat_i[6]
port 604 nsew
flabel metal2 s 38354 -960 38466 480 0 FreeSans 560 90 0 0 wbs_dat_i[7]
port 605 nsew
flabel metal2 s 41850 -960 41962 480 0 FreeSans 560 90 0 0 wbs_dat_i[8]
port 606 nsew
flabel metal2 s 45438 -960 45550 480 0 FreeSans 560 90 0 0 wbs_dat_i[9]
port 607 nsew
flabel metal2 s 9926 -960 10038 480 0 FreeSans 560 90 0 0 wbs_dat_o[0]
port 608 nsew
flabel metal2 s 50130 -960 50242 480 0 FreeSans 560 90 0 0 wbs_dat_o[10]
port 609 nsew
flabel metal2 s 53718 -960 53830 480 0 FreeSans 560 90 0 0 wbs_dat_o[11]
port 610 nsew
flabel metal2 s 57214 -960 57326 480 0 FreeSans 560 90 0 0 wbs_dat_o[12]
port 611 nsew
flabel metal2 s 60802 -960 60914 480 0 FreeSans 560 90 0 0 wbs_dat_o[13]
port 612 nsew
flabel metal2 s 64298 -960 64410 480 0 FreeSans 560 90 0 0 wbs_dat_o[14]
port 613 nsew
flabel metal2 s 67886 -960 67998 480 0 FreeSans 560 90 0 0 wbs_dat_o[15]
port 614 nsew
flabel metal2 s 71474 -960 71586 480 0 FreeSans 560 90 0 0 wbs_dat_o[16]
port 615 nsew
flabel metal2 s 74970 -960 75082 480 0 FreeSans 560 90 0 0 wbs_dat_o[17]
port 616 nsew
flabel metal2 s 78558 -960 78670 480 0 FreeSans 560 90 0 0 wbs_dat_o[18]
port 617 nsew
flabel metal2 s 82054 -960 82166 480 0 FreeSans 560 90 0 0 wbs_dat_o[19]
port 618 nsew
flabel metal2 s 14710 -960 14822 480 0 FreeSans 560 90 0 0 wbs_dat_o[1]
port 619 nsew
flabel metal2 s 85642 -960 85754 480 0 FreeSans 560 90 0 0 wbs_dat_o[20]
port 620 nsew
flabel metal2 s 89138 -960 89250 480 0 FreeSans 560 90 0 0 wbs_dat_o[21]
port 621 nsew
flabel metal2 s 92726 -960 92838 480 0 FreeSans 560 90 0 0 wbs_dat_o[22]
port 622 nsew
flabel metal2 s 96222 -960 96334 480 0 FreeSans 560 90 0 0 wbs_dat_o[23]
port 623 nsew
flabel metal2 s 99810 -960 99922 480 0 FreeSans 560 90 0 0 wbs_dat_o[24]
port 624 nsew
flabel metal2 s 103306 -960 103418 480 0 FreeSans 560 90 0 0 wbs_dat_o[25]
port 625 nsew
flabel metal2 s 106894 -960 107006 480 0 FreeSans 560 90 0 0 wbs_dat_o[26]
port 626 nsew
flabel metal2 s 110482 -960 110594 480 0 FreeSans 560 90 0 0 wbs_dat_o[27]
port 627 nsew
flabel metal2 s 113978 -960 114090 480 0 FreeSans 560 90 0 0 wbs_dat_o[28]
port 628 nsew
flabel metal2 s 117566 -960 117678 480 0 FreeSans 560 90 0 0 wbs_dat_o[29]
port 629 nsew
flabel metal2 s 19402 -960 19514 480 0 FreeSans 560 90 0 0 wbs_dat_o[2]
port 630 nsew
flabel metal2 s 121062 -960 121174 480 0 FreeSans 560 90 0 0 wbs_dat_o[30]
port 631 nsew
flabel metal2 s 124650 -960 124762 480 0 FreeSans 560 90 0 0 wbs_dat_o[31]
port 632 nsew
flabel metal2 s 24186 -960 24298 480 0 FreeSans 560 90 0 0 wbs_dat_o[3]
port 633 nsew
flabel metal2 s 28878 -960 28990 480 0 FreeSans 560 90 0 0 wbs_dat_o[4]
port 634 nsew
flabel metal2 s 32374 -960 32486 480 0 FreeSans 560 90 0 0 wbs_dat_o[5]
port 635 nsew
flabel metal2 s 35962 -960 36074 480 0 FreeSans 560 90 0 0 wbs_dat_o[6]
port 636 nsew
flabel metal2 s 39550 -960 39662 480 0 FreeSans 560 90 0 0 wbs_dat_o[7]
port 637 nsew
flabel metal2 s 43046 -960 43158 480 0 FreeSans 560 90 0 0 wbs_dat_o[8]
port 638 nsew
flabel metal2 s 46634 -960 46746 480 0 FreeSans 560 90 0 0 wbs_dat_o[9]
port 639 nsew
flabel metal2 s 11122 -960 11234 480 0 FreeSans 560 90 0 0 wbs_sel_i[0]
port 640 nsew
flabel metal2 s 15906 -960 16018 480 0 FreeSans 560 90 0 0 wbs_sel_i[1]
port 641 nsew
flabel metal2 s 20598 -960 20710 480 0 FreeSans 560 90 0 0 wbs_sel_i[2]
port 642 nsew
flabel metal2 s 25290 -960 25402 480 0 FreeSans 560 90 0 0 wbs_sel_i[3]
port 643 nsew
flabel metal2 s 5234 -960 5346 480 0 FreeSans 560 90 0 0 wbs_stb_i
port 644 nsew
flabel metal2 s 6430 -960 6542 480 0 FreeSans 560 90 0 0 wbs_we_i
port 645 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
